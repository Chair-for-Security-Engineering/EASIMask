// Generator : SpinalHDL v1.6.2    git head : e20135930d099f5d7469bbea4f2ca5d14698f642
// Component : G4MulTIMaskedN
// Git hash  : e20135930d099f5d7469bbea4f2ca5d14698f642

`timescale 1ns/1ps 

module G4MulTIMaskedN (
  input      [1:0]    io_x_0,
  input      [1:0]    io_x_1,
  input      [1:0]    io_x_2,
  input      [1:0]    io_x_3,
  input      [1:0]    io_x_4,
  input      [1:0]    io_x_5,
  input      [1:0]    io_x_6,
  input      [1:0]    io_x_7,
  input      [1:0]    io_x_8,
  input      [1:0]    io_y_0,
  input      [1:0]    io_y_1,
  input      [1:0]    io_y_2,
  input      [1:0]    io_y_3,
  input      [1:0]    io_y_4,
  input      [1:0]    io_y_5,
  input      [1:0]    io_y_6,
  input      [1:0]    io_y_7,
  input      [1:0]    io_y_8,
  output     [1:0]    io_z_0,
  output     [1:0]    io_z_1,
  output     [1:0]    io_z_2,
  output     [1:0]    io_z_3,
  output     [1:0]    io_z_4,
  output     [1:0]    io_z_5,
  output     [1:0]    io_z_6,
  output     [1:0]    io_z_7,
  output     [1:0]    io_z_8,
  input               clk,
  input               reset
);

  wire                dummy;
  wire                a_0;
  wire                a_1;
  wire                a_2;
  wire                a_3;
  wire                a_4;
  wire                a_5;
  wire                a_6;
  wire                a_7;
  wire                a_8;
  wire                b_0;
  wire                b_1;
  wire                b_2;
  wire                b_3;
  wire                b_4;
  wire                b_5;
  wire                b_6;
  wire                b_7;
  wire                b_8;
  wire                c_0;
  wire                c_1;
  wire                c_2;
  wire                c_3;
  wire                c_4;
  wire                c_5;
  wire                c_6;
  wire                c_7;
  wire                c_8;
  wire                d_0;
  wire                d_1;
  wire                d_2;
  wire                d_3;
  wire                d_4;
  wire                d_5;
  wire                d_6;
  wire                d_7;
  wire                d_8;
  reg        [8:0]    e_0;
  reg        [8:0]    e_1;
  reg        [8:0]    e_2;
  reg        [8:0]    e_3;
  reg        [8:0]    e_4;
  reg        [8:0]    e_5;
  reg        [8:0]    e_6;
  reg        [8:0]    e_7;
  reg        [8:0]    e_8;
  reg        [8:0]    f_0;
  reg        [8:0]    f_1;
  reg        [8:0]    f_2;
  reg        [8:0]    f_3;
  reg        [8:0]    f_4;
  reg        [8:0]    f_5;
  reg        [8:0]    f_6;
  reg        [8:0]    f_7;
  reg        [8:0]    f_8;
  wire                ac_0;
  wire                ac_1;
  wire                ac_2;
  wire                ac_3;
  wire                ac_4;
  wire                ac_5;
  wire                ac_6;
  wire                ac_7;
  wire                ac_8;
  wire                ac_9;
  wire                ac_10;
  wire                ac_11;
  wire                ac_12;
  wire                ac_13;
  wire                ac_14;
  wire                ac_15;
  wire                ac_16;
  wire                ac_17;
  wire                ac_18;
  wire                ac_19;
  wire                ac_20;
  wire                ac_21;
  wire                ac_22;
  wire                ac_23;
  wire                ac_24;
  wire                ac_25;
  wire                ac_26;
  wire                ac_27;
  wire                ac_28;
  wire                ac_29;
  wire                ac_30;
  wire                ac_31;
  wire                ac_32;
  wire                ac_33;
  wire                ac_34;
  wire                ac_35;
  wire                ac_36;
  wire                ac_37;
  wire                ac_38;
  wire                ac_39;
  wire                ac_40;
  wire                ac_41;
  wire                ac_42;
  wire                ac_43;
  wire                ac_44;
  wire                ac_45;
  wire                ac_46;
  wire                ac_47;
  wire                ac_48;
  wire                ac_49;
  wire                ac_50;
  wire                ac_51;
  wire                ac_52;
  wire                ac_53;
  wire                ac_54;
  wire                ac_55;
  wire                ac_56;
  wire                ac_57;
  wire                ac_58;
  wire                ac_59;
  wire                ac_60;
  wire                ac_61;
  wire                ac_62;
  wire                ac_63;
  wire                ac_64;
  wire                ac_65;
  wire                ac_66;
  wire                ac_67;
  wire                ac_68;
  wire                ac_69;
  wire                ac_70;
  wire                ac_71;
  wire                ac_72;
  wire                ac_73;
  wire                ac_74;
  wire                ac_75;
  wire                ac_76;
  wire                ac_77;
  wire                ac_78;
  wire                ac_79;
  wire                ac_80;
  wire                ad_0;
  wire                ad_1;
  wire                ad_2;
  wire                ad_3;
  wire                ad_4;
  wire                ad_5;
  wire                ad_6;
  wire                ad_7;
  wire                ad_8;
  wire                ad_9;
  wire                ad_10;
  wire                ad_11;
  wire                ad_12;
  wire                ad_13;
  wire                ad_14;
  wire                ad_15;
  wire                ad_16;
  wire                ad_17;
  wire                ad_18;
  wire                ad_19;
  wire                ad_20;
  wire                ad_21;
  wire                ad_22;
  wire                ad_23;
  wire                ad_24;
  wire                ad_25;
  wire                ad_26;
  wire                ad_27;
  wire                ad_28;
  wire                ad_29;
  wire                ad_30;
  wire                ad_31;
  wire                ad_32;
  wire                ad_33;
  wire                ad_34;
  wire                ad_35;
  wire                ad_36;
  wire                ad_37;
  wire                ad_38;
  wire                ad_39;
  wire                ad_40;
  wire                ad_41;
  wire                ad_42;
  wire                ad_43;
  wire                ad_44;
  wire                ad_45;
  wire                ad_46;
  wire                ad_47;
  wire                ad_48;
  wire                ad_49;
  wire                ad_50;
  wire                ad_51;
  wire                ad_52;
  wire                ad_53;
  wire                ad_54;
  wire                ad_55;
  wire                ad_56;
  wire                ad_57;
  wire                ad_58;
  wire                ad_59;
  wire                ad_60;
  wire                ad_61;
  wire                ad_62;
  wire                ad_63;
  wire                ad_64;
  wire                ad_65;
  wire                ad_66;
  wire                ad_67;
  wire                ad_68;
  wire                ad_69;
  wire                ad_70;
  wire                ad_71;
  wire                ad_72;
  wire                ad_73;
  wire                ad_74;
  wire                ad_75;
  wire                ad_76;
  wire                ad_77;
  wire                ad_78;
  wire                ad_79;
  wire                ad_80;
  wire                bc_0;
  wire                bc_1;
  wire                bc_2;
  wire                bc_3;
  wire                bc_4;
  wire                bc_5;
  wire                bc_6;
  wire                bc_7;
  wire                bc_8;
  wire                bc_9;
  wire                bc_10;
  wire                bc_11;
  wire                bc_12;
  wire                bc_13;
  wire                bc_14;
  wire                bc_15;
  wire                bc_16;
  wire                bc_17;
  wire                bc_18;
  wire                bc_19;
  wire                bc_20;
  wire                bc_21;
  wire                bc_22;
  wire                bc_23;
  wire                bc_24;
  wire                bc_25;
  wire                bc_26;
  wire                bc_27;
  wire                bc_28;
  wire                bc_29;
  wire                bc_30;
  wire                bc_31;
  wire                bc_32;
  wire                bc_33;
  wire                bc_34;
  wire                bc_35;
  wire                bc_36;
  wire                bc_37;
  wire                bc_38;
  wire                bc_39;
  wire                bc_40;
  wire                bc_41;
  wire                bc_42;
  wire                bc_43;
  wire                bc_44;
  wire                bc_45;
  wire                bc_46;
  wire                bc_47;
  wire                bc_48;
  wire                bc_49;
  wire                bc_50;
  wire                bc_51;
  wire                bc_52;
  wire                bc_53;
  wire                bc_54;
  wire                bc_55;
  wire                bc_56;
  wire                bc_57;
  wire                bc_58;
  wire                bc_59;
  wire                bc_60;
  wire                bc_61;
  wire                bc_62;
  wire                bc_63;
  wire                bc_64;
  wire                bc_65;
  wire                bc_66;
  wire                bc_67;
  wire                bc_68;
  wire                bc_69;
  wire                bc_70;
  wire                bc_71;
  wire                bc_72;
  wire                bc_73;
  wire                bc_74;
  wire                bc_75;
  wire                bc_76;
  wire                bc_77;
  wire                bc_78;
  wire                bc_79;
  wire                bc_80;
  wire                bd_0;
  wire                bd_1;
  wire                bd_2;
  wire                bd_3;
  wire                bd_4;
  wire                bd_5;
  wire                bd_6;
  wire                bd_7;
  wire                bd_8;
  wire                bd_9;
  wire                bd_10;
  wire                bd_11;
  wire                bd_12;
  wire                bd_13;
  wire                bd_14;
  wire                bd_15;
  wire                bd_16;
  wire                bd_17;
  wire                bd_18;
  wire                bd_19;
  wire                bd_20;
  wire                bd_21;
  wire                bd_22;
  wire                bd_23;
  wire                bd_24;
  wire                bd_25;
  wire                bd_26;
  wire                bd_27;
  wire                bd_28;
  wire                bd_29;
  wire                bd_30;
  wire                bd_31;
  wire                bd_32;
  wire                bd_33;
  wire                bd_34;
  wire                bd_35;
  wire                bd_36;
  wire                bd_37;
  wire                bd_38;
  wire                bd_39;
  wire                bd_40;
  wire                bd_41;
  wire                bd_42;
  wire                bd_43;
  wire                bd_44;
  wire                bd_45;
  wire                bd_46;
  wire                bd_47;
  wire                bd_48;
  wire                bd_49;
  wire                bd_50;
  wire                bd_51;
  wire                bd_52;
  wire                bd_53;
  wire                bd_54;
  wire                bd_55;
  wire                bd_56;
  wire                bd_57;
  wire                bd_58;
  wire                bd_59;
  wire                bd_60;
  wire                bd_61;
  wire                bd_62;
  wire                bd_63;
  wire                bd_64;
  wire                bd_65;
  wire                bd_66;
  wire                bd_67;
  wire                bd_68;
  wire                bd_69;
  wire                bd_70;
  wire                bd_71;
  wire                bd_72;
  wire                bd_73;
  wire                bd_74;
  wire                bd_75;
  wire                bd_76;
  wire                bd_77;
  wire                bd_78;
  wire                bd_79;
  wire                bd_80;

  assign dummy = 1'b0;
  assign a_0 = io_x_0[1];
  assign b_0 = io_x_0[0];
  assign c_0 = io_y_0[1];
  assign d_0 = io_y_0[0];
  assign a_1 = io_x_1[1];
  assign b_1 = io_x_1[0];
  assign c_1 = io_y_1[1];
  assign d_1 = io_y_1[0];
  assign a_2 = io_x_2[1];
  assign b_2 = io_x_2[0];
  assign c_2 = io_y_2[1];
  assign d_2 = io_y_2[0];
  assign a_3 = io_x_3[1];
  assign b_3 = io_x_3[0];
  assign c_3 = io_y_3[1];
  assign d_3 = io_y_3[0];
  assign a_4 = io_x_4[1];
  assign b_4 = io_x_4[0];
  assign c_4 = io_y_4[1];
  assign d_4 = io_y_4[0];
  assign a_5 = io_x_5[1];
  assign b_5 = io_x_5[0];
  assign c_5 = io_y_5[1];
  assign d_5 = io_y_5[0];
  assign a_6 = io_x_6[1];
  assign b_6 = io_x_6[0];
  assign c_6 = io_y_6[1];
  assign d_6 = io_y_6[0];
  assign a_7 = io_x_7[1];
  assign b_7 = io_x_7[0];
  assign c_7 = io_y_7[1];
  assign d_7 = io_y_7[0];
  assign a_8 = io_x_8[1];
  assign b_8 = io_x_8[0];
  assign c_8 = io_y_8[1];
  assign d_8 = io_y_8[0];
  assign ac_0 = (a_0 && c_0);
  assign ad_0 = (a_0 && d_0);
  assign bc_0 = (b_0 && c_0);
  assign bd_0 = (b_0 && d_0);
  assign ac_1 = (a_0 && c_1);
  assign ad_1 = (a_0 && d_1);
  assign bc_1 = (b_0 && c_1);
  assign bd_1 = (b_0 && d_1);
  assign ac_2 = (a_0 && c_2);
  assign ad_2 = (a_0 && d_2);
  assign bc_2 = (b_0 && c_2);
  assign bd_2 = (b_0 && d_2);
  assign ac_3 = (a_0 && c_3);
  assign ad_3 = (a_0 && d_3);
  assign bc_3 = (b_0 && c_3);
  assign bd_3 = (b_0 && d_3);
  assign ac_4 = (a_0 && c_4);
  assign ad_4 = (a_0 && d_4);
  assign bc_4 = (b_0 && c_4);
  assign bd_4 = (b_0 && d_4);
  assign ac_5 = (a_0 && c_5);
  assign ad_5 = (a_0 && d_5);
  assign bc_5 = (b_0 && c_5);
  assign bd_5 = (b_0 && d_5);
  assign ac_6 = (a_0 && c_6);
  assign ad_6 = (a_0 && d_6);
  assign bc_6 = (b_0 && c_6);
  assign bd_6 = (b_0 && d_6);
  assign ac_7 = (a_0 && c_7);
  assign ad_7 = (a_0 && d_7);
  assign bc_7 = (b_0 && c_7);
  assign bd_7 = (b_0 && d_7);
  assign ac_8 = (a_0 && c_8);
  assign ad_8 = (a_0 && d_8);
  assign bc_8 = (b_0 && c_8);
  assign bd_8 = (b_0 && d_8);
  assign ac_9 = (a_1 && c_0);
  assign ad_9 = (a_1 && d_0);
  assign bc_9 = (b_1 && c_0);
  assign bd_9 = (b_1 && d_0);
  assign ac_10 = (a_1 && c_1);
  assign ad_10 = (a_1 && d_1);
  assign bc_10 = (b_1 && c_1);
  assign bd_10 = (b_1 && d_1);
  assign ac_11 = (a_1 && c_2);
  assign ad_11 = (a_1 && d_2);
  assign bc_11 = (b_1 && c_2);
  assign bd_11 = (b_1 && d_2);
  assign ac_12 = (a_1 && c_3);
  assign ad_12 = (a_1 && d_3);
  assign bc_12 = (b_1 && c_3);
  assign bd_12 = (b_1 && d_3);
  assign ac_13 = (a_1 && c_4);
  assign ad_13 = (a_1 && d_4);
  assign bc_13 = (b_1 && c_4);
  assign bd_13 = (b_1 && d_4);
  assign ac_14 = (a_1 && c_5);
  assign ad_14 = (a_1 && d_5);
  assign bc_14 = (b_1 && c_5);
  assign bd_14 = (b_1 && d_5);
  assign ac_15 = (a_1 && c_6);
  assign ad_15 = (a_1 && d_6);
  assign bc_15 = (b_1 && c_6);
  assign bd_15 = (b_1 && d_6);
  assign ac_16 = (a_1 && c_7);
  assign ad_16 = (a_1 && d_7);
  assign bc_16 = (b_1 && c_7);
  assign bd_16 = (b_1 && d_7);
  assign ac_17 = (a_1 && c_8);
  assign ad_17 = (a_1 && d_8);
  assign bc_17 = (b_1 && c_8);
  assign bd_17 = (b_1 && d_8);
  assign ac_18 = (a_2 && c_0);
  assign ad_18 = (a_2 && d_0);
  assign bc_18 = (b_2 && c_0);
  assign bd_18 = (b_2 && d_0);
  assign ac_19 = (a_2 && c_1);
  assign ad_19 = (a_2 && d_1);
  assign bc_19 = (b_2 && c_1);
  assign bd_19 = (b_2 && d_1);
  assign ac_20 = (a_2 && c_2);
  assign ad_20 = (a_2 && d_2);
  assign bc_20 = (b_2 && c_2);
  assign bd_20 = (b_2 && d_2);
  assign ac_21 = (a_2 && c_3);
  assign ad_21 = (a_2 && d_3);
  assign bc_21 = (b_2 && c_3);
  assign bd_21 = (b_2 && d_3);
  assign ac_22 = (a_2 && c_4);
  assign ad_22 = (a_2 && d_4);
  assign bc_22 = (b_2 && c_4);
  assign bd_22 = (b_2 && d_4);
  assign ac_23 = (a_2 && c_5);
  assign ad_23 = (a_2 && d_5);
  assign bc_23 = (b_2 && c_5);
  assign bd_23 = (b_2 && d_5);
  assign ac_24 = (a_2 && c_6);
  assign ad_24 = (a_2 && d_6);
  assign bc_24 = (b_2 && c_6);
  assign bd_24 = (b_2 && d_6);
  assign ac_25 = (a_2 && c_7);
  assign ad_25 = (a_2 && d_7);
  assign bc_25 = (b_2 && c_7);
  assign bd_25 = (b_2 && d_7);
  assign ac_26 = (a_2 && c_8);
  assign ad_26 = (a_2 && d_8);
  assign bc_26 = (b_2 && c_8);
  assign bd_26 = (b_2 && d_8);
  assign ac_27 = (a_3 && c_0);
  assign ad_27 = (a_3 && d_0);
  assign bc_27 = (b_3 && c_0);
  assign bd_27 = (b_3 && d_0);
  assign ac_28 = (a_3 && c_1);
  assign ad_28 = (a_3 && d_1);
  assign bc_28 = (b_3 && c_1);
  assign bd_28 = (b_3 && d_1);
  assign ac_29 = (a_3 && c_2);
  assign ad_29 = (a_3 && d_2);
  assign bc_29 = (b_3 && c_2);
  assign bd_29 = (b_3 && d_2);
  assign ac_30 = (a_3 && c_3);
  assign ad_30 = (a_3 && d_3);
  assign bc_30 = (b_3 && c_3);
  assign bd_30 = (b_3 && d_3);
  assign ac_31 = (a_3 && c_4);
  assign ad_31 = (a_3 && d_4);
  assign bc_31 = (b_3 && c_4);
  assign bd_31 = (b_3 && d_4);
  assign ac_32 = (a_3 && c_5);
  assign ad_32 = (a_3 && d_5);
  assign bc_32 = (b_3 && c_5);
  assign bd_32 = (b_3 && d_5);
  assign ac_33 = (a_3 && c_6);
  assign ad_33 = (a_3 && d_6);
  assign bc_33 = (b_3 && c_6);
  assign bd_33 = (b_3 && d_6);
  assign ac_34 = (a_3 && c_7);
  assign ad_34 = (a_3 && d_7);
  assign bc_34 = (b_3 && c_7);
  assign bd_34 = (b_3 && d_7);
  assign ac_35 = (a_3 && c_8);
  assign ad_35 = (a_3 && d_8);
  assign bc_35 = (b_3 && c_8);
  assign bd_35 = (b_3 && d_8);
  assign ac_36 = (a_4 && c_0);
  assign ad_36 = (a_4 && d_0);
  assign bc_36 = (b_4 && c_0);
  assign bd_36 = (b_4 && d_0);
  assign ac_37 = (a_4 && c_1);
  assign ad_37 = (a_4 && d_1);
  assign bc_37 = (b_4 && c_1);
  assign bd_37 = (b_4 && d_1);
  assign ac_38 = (a_4 && c_2);
  assign ad_38 = (a_4 && d_2);
  assign bc_38 = (b_4 && c_2);
  assign bd_38 = (b_4 && d_2);
  assign ac_39 = (a_4 && c_3);
  assign ad_39 = (a_4 && d_3);
  assign bc_39 = (b_4 && c_3);
  assign bd_39 = (b_4 && d_3);
  assign ac_40 = (a_4 && c_4);
  assign ad_40 = (a_4 && d_4);
  assign bc_40 = (b_4 && c_4);
  assign bd_40 = (b_4 && d_4);
  assign ac_41 = (a_4 && c_5);
  assign ad_41 = (a_4 && d_5);
  assign bc_41 = (b_4 && c_5);
  assign bd_41 = (b_4 && d_5);
  assign ac_42 = (a_4 && c_6);
  assign ad_42 = (a_4 && d_6);
  assign bc_42 = (b_4 && c_6);
  assign bd_42 = (b_4 && d_6);
  assign ac_43 = (a_4 && c_7);
  assign ad_43 = (a_4 && d_7);
  assign bc_43 = (b_4 && c_7);
  assign bd_43 = (b_4 && d_7);
  assign ac_44 = (a_4 && c_8);
  assign ad_44 = (a_4 && d_8);
  assign bc_44 = (b_4 && c_8);
  assign bd_44 = (b_4 && d_8);
  assign ac_45 = (a_5 && c_0);
  assign ad_45 = (a_5 && d_0);
  assign bc_45 = (b_5 && c_0);
  assign bd_45 = (b_5 && d_0);
  assign ac_46 = (a_5 && c_1);
  assign ad_46 = (a_5 && d_1);
  assign bc_46 = (b_5 && c_1);
  assign bd_46 = (b_5 && d_1);
  assign ac_47 = (a_5 && c_2);
  assign ad_47 = (a_5 && d_2);
  assign bc_47 = (b_5 && c_2);
  assign bd_47 = (b_5 && d_2);
  assign ac_48 = (a_5 && c_3);
  assign ad_48 = (a_5 && d_3);
  assign bc_48 = (b_5 && c_3);
  assign bd_48 = (b_5 && d_3);
  assign ac_49 = (a_5 && c_4);
  assign ad_49 = (a_5 && d_4);
  assign bc_49 = (b_5 && c_4);
  assign bd_49 = (b_5 && d_4);
  assign ac_50 = (a_5 && c_5);
  assign ad_50 = (a_5 && d_5);
  assign bc_50 = (b_5 && c_5);
  assign bd_50 = (b_5 && d_5);
  assign ac_51 = (a_5 && c_6);
  assign ad_51 = (a_5 && d_6);
  assign bc_51 = (b_5 && c_6);
  assign bd_51 = (b_5 && d_6);
  assign ac_52 = (a_5 && c_7);
  assign ad_52 = (a_5 && d_7);
  assign bc_52 = (b_5 && c_7);
  assign bd_52 = (b_5 && d_7);
  assign ac_53 = (a_5 && c_8);
  assign ad_53 = (a_5 && d_8);
  assign bc_53 = (b_5 && c_8);
  assign bd_53 = (b_5 && d_8);
  assign ac_54 = (a_6 && c_0);
  assign ad_54 = (a_6 && d_0);
  assign bc_54 = (b_6 && c_0);
  assign bd_54 = (b_6 && d_0);
  assign ac_55 = (a_6 && c_1);
  assign ad_55 = (a_6 && d_1);
  assign bc_55 = (b_6 && c_1);
  assign bd_55 = (b_6 && d_1);
  assign ac_56 = (a_6 && c_2);
  assign ad_56 = (a_6 && d_2);
  assign bc_56 = (b_6 && c_2);
  assign bd_56 = (b_6 && d_2);
  assign ac_57 = (a_6 && c_3);
  assign ad_57 = (a_6 && d_3);
  assign bc_57 = (b_6 && c_3);
  assign bd_57 = (b_6 && d_3);
  assign ac_58 = (a_6 && c_4);
  assign ad_58 = (a_6 && d_4);
  assign bc_58 = (b_6 && c_4);
  assign bd_58 = (b_6 && d_4);
  assign ac_59 = (a_6 && c_5);
  assign ad_59 = (a_6 && d_5);
  assign bc_59 = (b_6 && c_5);
  assign bd_59 = (b_6 && d_5);
  assign ac_60 = (a_6 && c_6);
  assign ad_60 = (a_6 && d_6);
  assign bc_60 = (b_6 && c_6);
  assign bd_60 = (b_6 && d_6);
  assign ac_61 = (a_6 && c_7);
  assign ad_61 = (a_6 && d_7);
  assign bc_61 = (b_6 && c_7);
  assign bd_61 = (b_6 && d_7);
  assign ac_62 = (a_6 && c_8);
  assign ad_62 = (a_6 && d_8);
  assign bc_62 = (b_6 && c_8);
  assign bd_62 = (b_6 && d_8);
  assign ac_63 = (a_7 && c_0);
  assign ad_63 = (a_7 && d_0);
  assign bc_63 = (b_7 && c_0);
  assign bd_63 = (b_7 && d_0);
  assign ac_64 = (a_7 && c_1);
  assign ad_64 = (a_7 && d_1);
  assign bc_64 = (b_7 && c_1);
  assign bd_64 = (b_7 && d_1);
  assign ac_65 = (a_7 && c_2);
  assign ad_65 = (a_7 && d_2);
  assign bc_65 = (b_7 && c_2);
  assign bd_65 = (b_7 && d_2);
  assign ac_66 = (a_7 && c_3);
  assign ad_66 = (a_7 && d_3);
  assign bc_66 = (b_7 && c_3);
  assign bd_66 = (b_7 && d_3);
  assign ac_67 = (a_7 && c_4);
  assign ad_67 = (a_7 && d_4);
  assign bc_67 = (b_7 && c_4);
  assign bd_67 = (b_7 && d_4);
  assign ac_68 = (a_7 && c_5);
  assign ad_68 = (a_7 && d_5);
  assign bc_68 = (b_7 && c_5);
  assign bd_68 = (b_7 && d_5);
  assign ac_69 = (a_7 && c_6);
  assign ad_69 = (a_7 && d_6);
  assign bc_69 = (b_7 && c_6);
  assign bd_69 = (b_7 && d_6);
  assign ac_70 = (a_7 && c_7);
  assign ad_70 = (a_7 && d_7);
  assign bc_70 = (b_7 && c_7);
  assign bd_70 = (b_7 && d_7);
  assign ac_71 = (a_7 && c_8);
  assign ad_71 = (a_7 && d_8);
  assign bc_71 = (b_7 && c_8);
  assign bd_71 = (b_7 && d_8);
  assign ac_72 = (a_8 && c_0);
  assign ad_72 = (a_8 && d_0);
  assign bc_72 = (b_8 && c_0);
  assign bd_72 = (b_8 && d_0);
  assign ac_73 = (a_8 && c_1);
  assign ad_73 = (a_8 && d_1);
  assign bc_73 = (b_8 && c_1);
  assign bd_73 = (b_8 && d_1);
  assign ac_74 = (a_8 && c_2);
  assign ad_74 = (a_8 && d_2);
  assign bc_74 = (b_8 && c_2);
  assign bd_74 = (b_8 && d_2);
  assign ac_75 = (a_8 && c_3);
  assign ad_75 = (a_8 && d_3);
  assign bc_75 = (b_8 && c_3);
  assign bd_75 = (b_8 && d_3);
  assign ac_76 = (a_8 && c_4);
  assign ad_76 = (a_8 && d_4);
  assign bc_76 = (b_8 && c_4);
  assign bd_76 = (b_8 && d_4);
  assign ac_77 = (a_8 && c_5);
  assign ad_77 = (a_8 && d_5);
  assign bc_77 = (b_8 && c_5);
  assign bd_77 = (b_8 && d_5);
  assign ac_78 = (a_8 && c_6);
  assign ad_78 = (a_8 && d_6);
  assign bc_78 = (b_8 && c_6);
  assign bd_78 = (b_8 && d_6);
  assign ac_79 = (a_8 && c_7);
  assign ad_79 = (a_8 && d_7);
  assign bc_79 = (b_8 && c_7);
  assign bd_79 = (b_8 && d_7);
  assign ac_80 = (a_8 && c_8);
  assign ad_80 = (a_8 && d_8);
  assign bc_80 = (b_8 && c_8);
  assign bd_80 = (b_8 && d_8);
  always @(*) begin
    e_0[8] = ((bc_0 ^ ad_0) ^ bd_0);
    e_0[0] = ((bc_10 ^ ad_10) ^ bd_10);
    e_0[1] = ((bc_20 ^ ad_20) ^ bd_20);
    e_0[2] = ((bc_30 ^ ad_30) ^ bd_30);
    e_0[3] = ((bc_40 ^ ad_40) ^ bd_40);
    e_0[4] = ((bc_50 ^ ad_50) ^ bd_50);
    e_0[5] = ((bc_60 ^ ad_60) ^ bd_60);
    e_0[6] = ((bc_70 ^ ad_70) ^ bd_70);
    e_0[7] = ((bc_80 ^ ad_80) ^ bd_80);
  end

  always @(*) begin
    f_0[8] = ((bc_0 ^ ad_0) ^ ac_0);
    f_0[0] = ((bc_10 ^ ad_10) ^ ac_10);
    f_0[1] = ((bc_20 ^ ad_20) ^ ac_20);
    f_0[2] = ((bc_30 ^ ad_30) ^ ac_30);
    f_0[3] = ((bc_40 ^ ad_40) ^ ac_40);
    f_0[4] = ((bc_50 ^ ad_50) ^ ac_50);
    f_0[5] = ((bc_60 ^ ad_60) ^ ac_60);
    f_0[6] = ((bc_70 ^ ad_70) ^ ac_70);
    f_0[7] = ((bc_80 ^ ad_80) ^ ac_80);
  end

  always @(*) begin
    e_1[0] = (((e_0[0] ^ bc_11) ^ ad_11) ^ bd_11);
    e_1[1] = (((e_0[1] ^ bc_2) ^ ad_2) ^ bd_2);
    e_1[2] = (((e_0[2] ^ bc_1) ^ ad_1) ^ bd_1);
    e_1[3] = (((e_0[3] ^ bc_4) ^ ad_4) ^ bd_4);
    e_1[4] = (((e_0[4] ^ bc_3) ^ ad_3) ^ bd_3);
    e_1[5] = (((e_0[5] ^ bc_6) ^ ad_6) ^ bd_6);
    e_1[6] = (((e_0[6] ^ bc_5) ^ ad_5) ^ bd_5);
    e_1[7] = (((e_0[7] ^ bc_8) ^ ad_8) ^ bd_8);
    e_1[8] = (((e_0[8] ^ bc_7) ^ ad_7) ^ bd_7);
  end

  always @(*) begin
    f_1[0] = (((f_0[0] ^ bc_11) ^ ad_11) ^ ac_11);
    f_1[1] = (((f_0[1] ^ bc_2) ^ ad_2) ^ ac_2);
    f_1[2] = (((f_0[2] ^ bc_1) ^ ad_1) ^ ac_1);
    f_1[3] = (((f_0[3] ^ bc_4) ^ ad_4) ^ ac_4);
    f_1[4] = (((f_0[4] ^ bc_3) ^ ad_3) ^ ac_3);
    f_1[5] = (((f_0[5] ^ bc_6) ^ ad_6) ^ ac_6);
    f_1[6] = (((f_0[6] ^ bc_5) ^ ad_5) ^ ac_5);
    f_1[7] = (((f_0[7] ^ bc_8) ^ ad_8) ^ ac_8);
    f_1[8] = (((f_0[8] ^ bc_7) ^ ad_7) ^ ac_7);
  end

  always @(*) begin
    e_2[0] = (((e_1[0] ^ bc_19) ^ ad_19) ^ bd_19);
    e_2[1] = (((e_1[1] ^ bc_18) ^ ad_18) ^ bd_18);
    e_2[2] = (((e_1[2] ^ bc_9) ^ ad_9) ^ bd_9);
    e_2[3] = (((e_1[3] ^ bc_13) ^ ad_13) ^ bd_13);
    e_2[4] = (((e_1[4] ^ bc_12) ^ ad_12) ^ bd_12);
    e_2[5] = (((e_1[5] ^ bc_15) ^ ad_15) ^ bd_15);
    e_2[6] = (((e_1[6] ^ bc_14) ^ ad_14) ^ bd_14);
    e_2[7] = (((e_1[7] ^ bc_17) ^ ad_17) ^ bd_17);
    e_2[8] = (((e_1[8] ^ bc_16) ^ ad_16) ^ bd_16);
  end

  always @(*) begin
    f_2[0] = (((f_1[0] ^ bc_19) ^ ad_19) ^ ac_19);
    f_2[1] = (((f_1[1] ^ bc_18) ^ ad_18) ^ ac_18);
    f_2[2] = (((f_1[2] ^ bc_9) ^ ad_9) ^ ac_9);
    f_2[3] = (((f_1[3] ^ bc_13) ^ ad_13) ^ ac_13);
    f_2[4] = (((f_1[4] ^ bc_12) ^ ad_12) ^ ac_12);
    f_2[5] = (((f_1[5] ^ bc_15) ^ ad_15) ^ ac_15);
    f_2[6] = (((f_1[6] ^ bc_14) ^ ad_14) ^ ac_14);
    f_2[7] = (((f_1[7] ^ bc_17) ^ ad_17) ^ ac_17);
    f_2[8] = (((f_1[8] ^ bc_16) ^ ad_16) ^ ac_16);
  end

  always @(*) begin
    e_3[0] = (((e_2[0] ^ bc_28) ^ ad_28) ^ bd_28);
    e_3[1] = (((e_2[1] ^ bc_27) ^ ad_27) ^ bd_27);
    e_3[2] = (((e_2[2] ^ bc_31) ^ ad_31) ^ bd_31);
    e_3[3] = (((e_2[3] ^ bc_22) ^ ad_22) ^ bd_22);
    e_3[4] = (((e_2[4] ^ bc_21) ^ ad_21) ^ bd_21);
    e_3[5] = (((e_2[5] ^ bc_24) ^ ad_24) ^ bd_24);
    e_3[6] = (((e_2[6] ^ bc_23) ^ ad_23) ^ bd_23);
    e_3[7] = (((e_2[7] ^ bc_26) ^ ad_26) ^ bd_26);
    e_3[8] = (((e_2[8] ^ bc_25) ^ ad_25) ^ bd_25);
  end

  always @(*) begin
    f_3[0] = (((f_2[0] ^ bc_28) ^ ad_28) ^ ac_28);
    f_3[1] = (((f_2[1] ^ bc_27) ^ ad_27) ^ ac_27);
    f_3[2] = (((f_2[2] ^ bc_31) ^ ad_31) ^ ac_31);
    f_3[3] = (((f_2[3] ^ bc_22) ^ ad_22) ^ ac_22);
    f_3[4] = (((f_2[4] ^ bc_21) ^ ad_21) ^ ac_21);
    f_3[5] = (((f_2[5] ^ bc_24) ^ ad_24) ^ ac_24);
    f_3[6] = (((f_2[6] ^ bc_23) ^ ad_23) ^ ac_23);
    f_3[7] = (((f_2[7] ^ bc_26) ^ ad_26) ^ ac_26);
    f_3[8] = (((f_2[8] ^ bc_25) ^ ad_25) ^ ac_25);
  end

  always @(*) begin
    e_4[0] = (((e_3[0] ^ bc_37) ^ ad_37) ^ bd_37);
    e_4[1] = (((e_3[1] ^ bc_36) ^ ad_36) ^ bd_36);
    e_4[2] = (((e_3[2] ^ bc_39) ^ ad_39) ^ bd_39);
    e_4[3] = (((e_3[3] ^ bc_38) ^ ad_38) ^ bd_38);
    e_4[4] = (((e_3[4] ^ bc_29) ^ ad_29) ^ bd_29);
    e_4[5] = (((e_3[5] ^ bc_33) ^ ad_33) ^ bd_33);
    e_4[6] = (((e_3[6] ^ bc_32) ^ ad_32) ^ bd_32);
    e_4[7] = (((e_3[7] ^ bc_35) ^ ad_35) ^ bd_35);
    e_4[8] = (((e_3[8] ^ bc_34) ^ ad_34) ^ bd_34);
  end

  always @(*) begin
    f_4[0] = (((f_3[0] ^ bc_37) ^ ad_37) ^ ac_37);
    f_4[1] = (((f_3[1] ^ bc_36) ^ ad_36) ^ ac_36);
    f_4[2] = (((f_3[2] ^ bc_39) ^ ad_39) ^ ac_39);
    f_4[3] = (((f_3[3] ^ bc_38) ^ ad_38) ^ ac_38);
    f_4[4] = (((f_3[4] ^ bc_29) ^ ad_29) ^ ac_29);
    f_4[5] = (((f_3[5] ^ bc_33) ^ ad_33) ^ ac_33);
    f_4[6] = (((f_3[6] ^ bc_32) ^ ad_32) ^ ac_32);
    f_4[7] = (((f_3[7] ^ bc_35) ^ ad_35) ^ ac_35);
    f_4[8] = (((f_3[8] ^ bc_34) ^ ad_34) ^ ac_34);
  end

  always @(*) begin
    e_5[0] = (((e_4[0] ^ bc_46) ^ ad_46) ^ bd_46);
    e_5[1] = (((e_4[1] ^ bc_45) ^ ad_45) ^ bd_45);
    e_5[2] = (((e_4[2] ^ bc_48) ^ ad_48) ^ bd_48);
    e_5[3] = (((e_4[3] ^ bc_47) ^ ad_47) ^ bd_47);
    e_5[4] = (((e_4[4] ^ bc_51) ^ ad_51) ^ bd_51);
    e_5[5] = (((e_4[5] ^ bc_42) ^ ad_42) ^ bd_42);
    e_5[6] = (((e_4[6] ^ bc_41) ^ ad_41) ^ bd_41);
    e_5[7] = (((e_4[7] ^ bc_44) ^ ad_44) ^ bd_44);
    e_5[8] = (((e_4[8] ^ bc_43) ^ ad_43) ^ bd_43);
  end

  always @(*) begin
    f_5[0] = (((f_4[0] ^ bc_46) ^ ad_46) ^ ac_46);
    f_5[1] = (((f_4[1] ^ bc_45) ^ ad_45) ^ ac_45);
    f_5[2] = (((f_4[2] ^ bc_48) ^ ad_48) ^ ac_48);
    f_5[3] = (((f_4[3] ^ bc_47) ^ ad_47) ^ ac_47);
    f_5[4] = (((f_4[4] ^ bc_51) ^ ad_51) ^ ac_51);
    f_5[5] = (((f_4[5] ^ bc_42) ^ ad_42) ^ ac_42);
    f_5[6] = (((f_4[6] ^ bc_41) ^ ad_41) ^ ac_41);
    f_5[7] = (((f_4[7] ^ bc_44) ^ ad_44) ^ ac_44);
    f_5[8] = (((f_4[8] ^ bc_43) ^ ad_43) ^ ac_43);
  end

  always @(*) begin
    e_6[0] = (((e_5[0] ^ bc_55) ^ ad_55) ^ bd_55);
    e_6[1] = (((e_5[1] ^ bc_54) ^ ad_54) ^ bd_54);
    e_6[2] = (((e_5[2] ^ bc_57) ^ ad_57) ^ bd_57);
    e_6[3] = (((e_5[3] ^ bc_56) ^ ad_56) ^ bd_56);
    e_6[4] = (((e_5[4] ^ bc_59) ^ ad_59) ^ bd_59);
    e_6[5] = (((e_5[5] ^ bc_58) ^ ad_58) ^ bd_58);
    e_6[6] = (((e_5[6] ^ bc_49) ^ ad_49) ^ bd_49);
    e_6[7] = (((e_5[7] ^ bc_53) ^ ad_53) ^ bd_53);
    e_6[8] = (((e_5[8] ^ bc_52) ^ ad_52) ^ bd_52);
  end

  always @(*) begin
    f_6[0] = (((f_5[0] ^ bc_55) ^ ad_55) ^ ac_55);
    f_6[1] = (((f_5[1] ^ bc_54) ^ ad_54) ^ ac_54);
    f_6[2] = (((f_5[2] ^ bc_57) ^ ad_57) ^ ac_57);
    f_6[3] = (((f_5[3] ^ bc_56) ^ ad_56) ^ ac_56);
    f_6[4] = (((f_5[4] ^ bc_59) ^ ad_59) ^ ac_59);
    f_6[5] = (((f_5[5] ^ bc_58) ^ ad_58) ^ ac_58);
    f_6[6] = (((f_5[6] ^ bc_49) ^ ad_49) ^ ac_49);
    f_6[7] = (((f_5[7] ^ bc_53) ^ ad_53) ^ ac_53);
    f_6[8] = (((f_5[8] ^ bc_52) ^ ad_52) ^ ac_52);
  end

  always @(*) begin
    e_7[0] = (((e_6[0] ^ bc_64) ^ ad_64) ^ bd_64);
    e_7[1] = (((e_6[1] ^ bc_63) ^ ad_63) ^ bd_63);
    e_7[2] = (((e_6[2] ^ bc_66) ^ ad_66) ^ bd_66);
    e_7[3] = (((e_6[3] ^ bc_65) ^ ad_65) ^ bd_65);
    e_7[4] = (((e_6[4] ^ bc_68) ^ ad_68) ^ bd_68);
    e_7[5] = (((e_6[5] ^ bc_67) ^ ad_67) ^ bd_67);
    e_7[6] = (((e_6[6] ^ bc_71) ^ ad_71) ^ bd_71);
    e_7[7] = (((e_6[7] ^ bc_62) ^ ad_62) ^ bd_62);
    e_7[8] = (((e_6[8] ^ bc_61) ^ ad_61) ^ bd_61);
  end

  always @(*) begin
    f_7[0] = (((f_6[0] ^ bc_64) ^ ad_64) ^ ac_64);
    f_7[1] = (((f_6[1] ^ bc_63) ^ ad_63) ^ ac_63);
    f_7[2] = (((f_6[2] ^ bc_66) ^ ad_66) ^ ac_66);
    f_7[3] = (((f_6[3] ^ bc_65) ^ ad_65) ^ ac_65);
    f_7[4] = (((f_6[4] ^ bc_68) ^ ad_68) ^ ac_68);
    f_7[5] = (((f_6[5] ^ bc_67) ^ ad_67) ^ ac_67);
    f_7[6] = (((f_6[6] ^ bc_71) ^ ad_71) ^ ac_71);
    f_7[7] = (((f_6[7] ^ bc_62) ^ ad_62) ^ ac_62);
    f_7[8] = (((f_6[8] ^ bc_61) ^ ad_61) ^ ac_61);
  end

  always @(*) begin
    e_8[0] = (((e_7[0] ^ bc_73) ^ ad_73) ^ bd_73);
    e_8[1] = (((e_7[1] ^ bc_72) ^ ad_72) ^ bd_72);
    e_8[2] = (((e_7[2] ^ bc_75) ^ ad_75) ^ bd_75);
    e_8[3] = (((e_7[3] ^ bc_74) ^ ad_74) ^ bd_74);
    e_8[4] = (((e_7[4] ^ bc_77) ^ ad_77) ^ bd_77);
    e_8[5] = (((e_7[5] ^ bc_76) ^ ad_76) ^ bd_76);
    e_8[6] = (((e_7[6] ^ bc_79) ^ ad_79) ^ bd_79);
    e_8[7] = (((e_7[7] ^ bc_78) ^ ad_78) ^ bd_78);
    e_8[8] = (((e_7[8] ^ bc_69) ^ ad_69) ^ bd_69);
  end

  always @(*) begin
    f_8[0] = (((f_7[0] ^ bc_73) ^ ad_73) ^ ac_73);
    f_8[1] = (((f_7[1] ^ bc_72) ^ ad_72) ^ ac_72);
    f_8[2] = (((f_7[2] ^ bc_75) ^ ad_75) ^ ac_75);
    f_8[3] = (((f_7[3] ^ bc_74) ^ ad_74) ^ ac_74);
    f_8[4] = (((f_7[4] ^ bc_77) ^ ad_77) ^ ac_77);
    f_8[5] = (((f_7[5] ^ bc_76) ^ ad_76) ^ ac_76);
    f_8[6] = (((f_7[6] ^ bc_79) ^ ad_79) ^ ac_79);
    f_8[7] = (((f_7[7] ^ bc_78) ^ ad_78) ^ ac_78);
    f_8[8] = (((f_7[8] ^ bc_69) ^ ad_69) ^ ac_69);
  end

  assign io_z_0 = {e_8[0],f_8[0]};
  assign io_z_1 = {e_8[1],f_8[1]};
  assign io_z_2 = {e_8[2],f_8[2]};
  assign io_z_3 = {e_8[3],f_8[3]};
  assign io_z_4 = {e_8[4],f_8[4]};
  assign io_z_5 = {e_8[5],f_8[5]};
  assign io_z_6 = {e_8[6],f_8[6]};
  assign io_z_7 = {e_8[7],f_8[7]};
  assign io_z_8 = {e_8[8],f_8[8]};

endmodule
