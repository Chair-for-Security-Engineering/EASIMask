// Generator : SpinalHDL v1.6.2    git head : e20135930d099f5d7469bbea4f2ca5d14698f642
// Component : G256InvTIMaskedN
// Git hash  : e20135930d099f5d7469bbea4f2ca5d14698f642

`timescale 1ns/1ps 

module G256InvTIMaskedN (
  input      [7:0]    io_x_0,
  input      [7:0]    io_x_1,
  input      [7:0]    io_x_2,
  input      [7:0]    io_x_3,
  input      [7:0]    io_x_4,
  input      [7:0]    io_x_5,
  input      [7:0]    io_x_6,
  input      [7:0]    io_x_7,
  input      [7:0]    io_x_8,
  input      [7:0]    io_x_9,
  input      [7:0]    io_x_10,
  input      [7:0]    io_x_11,
  input      [7:0]    io_x_12,
  output     [7:0]    io_z_0,
  output     [7:0]    io_z_1,
  output     [7:0]    io_z_2,
  output     [7:0]    io_z_3,
  output     [7:0]    io_z_4,
  output     [7:0]    io_z_5,
  output     [7:0]    io_z_6,
  output     [7:0]    io_z_7,
  output     [7:0]    io_z_8,
  output     [7:0]    io_z_9,
  output     [7:0]    io_z_10,
  output     [7:0]    io_z_11,
  output     [7:0]    io_z_12,
  input               clk,
  input               reset
);

  wire       [3:0]    inv_io_x_0;
  wire       [3:0]    inv_io_x_1;
  wire       [3:0]    inv_io_x_2;
  wire       [3:0]    inv_io_x_3;
  wire       [3:0]    inv_io_x_4;
  wire       [3:0]    inv_io_x_5;
  wire       [3:0]    inv_io_x_6;
  wire       [3:0]    inv_io_x_7;
  wire       [3:0]    inv_io_x_8;
  wire       [3:0]    inv_io_x_9;
  wire       [3:0]    inv_io_x_10;
  wire       [3:0]    inv_io_x_11;
  wire       [3:0]    inv_io_x_12;
  wire       [3:0]    mul1_io_z_0;
  wire       [3:0]    mul1_io_z_1;
  wire       [3:0]    mul1_io_z_2;
  wire       [3:0]    mul1_io_z_3;
  wire       [3:0]    mul1_io_z_4;
  wire       [3:0]    mul1_io_z_5;
  wire       [3:0]    mul1_io_z_6;
  wire       [3:0]    mul1_io_z_7;
  wire       [3:0]    mul1_io_z_8;
  wire       [3:0]    mul1_io_z_9;
  wire       [3:0]    mul1_io_z_10;
  wire       [3:0]    mul1_io_z_11;
  wire       [3:0]    mul1_io_z_12;
  wire       [3:0]    mul2_io_z_0;
  wire       [3:0]    mul2_io_z_1;
  wire       [3:0]    mul2_io_z_2;
  wire       [3:0]    mul2_io_z_3;
  wire       [3:0]    mul2_io_z_4;
  wire       [3:0]    mul2_io_z_5;
  wire       [3:0]    mul2_io_z_6;
  wire       [3:0]    mul2_io_z_7;
  wire       [3:0]    mul2_io_z_8;
  wire       [3:0]    mul2_io_z_9;
  wire       [3:0]    mul2_io_z_10;
  wire       [3:0]    mul2_io_z_11;
  wire       [3:0]    mul2_io_z_12;
  wire       [3:0]    mul3_io_z_0;
  wire       [3:0]    mul3_io_z_1;
  wire       [3:0]    mul3_io_z_2;
  wire       [3:0]    mul3_io_z_3;
  wire       [3:0]    mul3_io_z_4;
  wire       [3:0]    mul3_io_z_5;
  wire       [3:0]    mul3_io_z_6;
  wire       [3:0]    mul3_io_z_7;
  wire       [3:0]    mul3_io_z_8;
  wire       [3:0]    mul3_io_z_9;
  wire       [3:0]    mul3_io_z_10;
  wire       [3:0]    mul3_io_z_11;
  wire       [3:0]    mul3_io_z_12;
  wire       [3:0]    inv_io_z_0;
  wire       [3:0]    inv_io_z_1;
  wire       [3:0]    inv_io_z_2;
  wire       [3:0]    inv_io_z_3;
  wire       [3:0]    inv_io_z_4;
  wire       [3:0]    inv_io_z_5;
  wire       [3:0]    inv_io_z_6;
  wire       [3:0]    inv_io_z_7;
  wire       [3:0]    inv_io_z_8;
  wire       [3:0]    inv_io_z_9;
  wire       [3:0]    inv_io_z_10;
  wire       [3:0]    inv_io_z_11;
  wire       [3:0]    inv_io_z_12;
  wire       [3:0]    g16SqSc_13_io_x;
  wire       [3:0]    g16SqSc_14_io_x;
  wire       [3:0]    g16SqSc_15_io_x;
  wire       [3:0]    g16SqSc_16_io_x;
  wire       [3:0]    g16SqSc_17_io_x;
  wire       [3:0]    g16SqSc_18_io_x;
  wire       [3:0]    g16SqSc_19_io_x;
  wire       [3:0]    g16SqSc_20_io_x;
  wire       [3:0]    g16SqSc_21_io_x;
  wire       [3:0]    g16SqSc_22_io_x;
  wire       [3:0]    g16SqSc_23_io_x;
  wire       [3:0]    g16SqSc_24_io_x;
  wire       [3:0]    g16SqSc_25_io_x;
  wire                dummy;
  wire       [3:0]    a_0;
  wire       [3:0]    a_1;
  wire       [3:0]    a_2;
  wire       [3:0]    a_3;
  wire       [3:0]    a_4;
  wire       [3:0]    a_5;
  wire       [3:0]    a_6;
  wire       [3:0]    a_7;
  wire       [3:0]    a_8;
  wire       [3:0]    a_9;
  wire       [3:0]    a_10;
  wire       [3:0]    a_11;
  wire       [3:0]    a_12;
  wire       [3:0]    b_0;
  wire       [3:0]    b_1;
  wire       [3:0]    b_2;
  wire       [3:0]    b_3;
  wire       [3:0]    b_4;
  wire       [3:0]    b_5;
  wire       [3:0]    b_6;
  wire       [3:0]    b_7;
  wire       [3:0]    b_8;
  wire       [3:0]    b_9;
  wire       [3:0]    b_10;
  wire       [3:0]    b_11;
  wire       [3:0]    b_12;
  wire       [3:0]    c_0;
  wire       [3:0]    c_1;
  wire       [3:0]    c_2;
  wire       [3:0]    c_3;
  wire       [3:0]    c_4;
  wire       [3:0]    c_5;
  wire       [3:0]    c_6;
  wire       [3:0]    c_7;
  wire       [3:0]    c_8;
  wire       [3:0]    c_9;
  wire       [3:0]    c_10;
  wire       [3:0]    c_11;
  wire       [3:0]    c_12;
  wire       [3:0]    d_0;
  wire       [3:0]    d_1;
  wire       [3:0]    d_2;
  wire       [3:0]    d_3;
  wire       [3:0]    d_4;
  wire       [3:0]    d_5;
  wire       [3:0]    d_6;
  wire       [3:0]    d_7;
  wire       [3:0]    d_8;
  wire       [3:0]    d_9;
  wire       [3:0]    d_10;
  wire       [3:0]    d_11;
  wire       [3:0]    d_12;
  wire       [3:0]    e_0;
  wire       [3:0]    e_1;
  wire       [3:0]    e_2;
  wire       [3:0]    e_3;
  wire       [3:0]    e_4;
  wire       [3:0]    e_5;
  wire       [3:0]    e_6;
  wire       [3:0]    e_7;
  wire       [3:0]    e_8;
  wire       [3:0]    e_9;
  wire       [3:0]    e_10;
  wire       [3:0]    e_11;
  wire       [3:0]    e_12;
  wire       [3:0]    f_0;
  wire       [3:0]    f_1;
  wire       [3:0]    f_2;
  wire       [3:0]    f_3;
  wire       [3:0]    f_4;
  wire       [3:0]    f_5;
  wire       [3:0]    f_6;
  wire       [3:0]    f_7;
  wire       [3:0]    f_8;
  wire       [3:0]    f_9;
  wire       [3:0]    f_10;
  wire       [3:0]    f_11;
  wire       [3:0]    f_12;
  wire       [3:0]    p_0;
  wire       [3:0]    p_1;
  wire       [3:0]    p_2;
  wire       [3:0]    p_3;
  wire       [3:0]    p_4;
  wire       [3:0]    p_5;
  wire       [3:0]    p_6;
  wire       [3:0]    p_7;
  wire       [3:0]    p_8;
  wire       [3:0]    p_9;
  wire       [3:0]    p_10;
  wire       [3:0]    p_11;
  wire       [3:0]    p_12;
  wire       [3:0]    q_0;
  wire       [3:0]    q_1;
  wire       [3:0]    q_2;
  wire       [3:0]    q_3;
  wire       [3:0]    q_4;
  wire       [3:0]    q_5;
  wire       [3:0]    q_6;
  wire       [3:0]    q_7;
  wire       [3:0]    q_8;
  wire       [3:0]    q_9;
  wire       [3:0]    q_10;
  wire       [3:0]    q_11;
  wire       [3:0]    q_12;

  G16MulTIMaskedN mul1 (
    .io_x_0     (a_0[3:0]           ), //i
    .io_x_1     (a_1[3:0]           ), //i
    .io_x_2     (a_2[3:0]           ), //i
    .io_x_3     (a_3[3:0]           ), //i
    .io_x_4     (a_4[3:0]           ), //i
    .io_x_5     (a_5[3:0]           ), //i
    .io_x_6     (a_6[3:0]           ), //i
    .io_x_7     (a_7[3:0]           ), //i
    .io_x_8     (a_8[3:0]           ), //i
    .io_x_9     (a_9[3:0]           ), //i
    .io_x_10    (a_10[3:0]          ), //i
    .io_x_11    (a_11[3:0]          ), //i
    .io_x_12    (a_12[3:0]          ), //i
    .io_y_0     (b_0[3:0]           ), //i
    .io_y_1     (b_1[3:0]           ), //i
    .io_y_2     (b_2[3:0]           ), //i
    .io_y_3     (b_3[3:0]           ), //i
    .io_y_4     (b_4[3:0]           ), //i
    .io_y_5     (b_5[3:0]           ), //i
    .io_y_6     (b_6[3:0]           ), //i
    .io_y_7     (b_7[3:0]           ), //i
    .io_y_8     (b_8[3:0]           ), //i
    .io_y_9     (b_9[3:0]           ), //i
    .io_y_10    (b_10[3:0]          ), //i
    .io_y_11    (b_11[3:0]          ), //i
    .io_y_12    (b_12[3:0]          ), //i
    .io_z_0     (mul1_io_z_0[3:0]   ), //o
    .io_z_1     (mul1_io_z_1[3:0]   ), //o
    .io_z_2     (mul1_io_z_2[3:0]   ), //o
    .io_z_3     (mul1_io_z_3[3:0]   ), //o
    .io_z_4     (mul1_io_z_4[3:0]   ), //o
    .io_z_5     (mul1_io_z_5[3:0]   ), //o
    .io_z_6     (mul1_io_z_6[3:0]   ), //o
    .io_z_7     (mul1_io_z_7[3:0]   ), //o
    .io_z_8     (mul1_io_z_8[3:0]   ), //o
    .io_z_9     (mul1_io_z_9[3:0]   ), //o
    .io_z_10    (mul1_io_z_10[3:0]  ), //o
    .io_z_11    (mul1_io_z_11[3:0]  ), //o
    .io_z_12    (mul1_io_z_12[3:0]  ), //o
    .clk        (clk                ), //i
    .reset      (reset              )  //i
  );
  G16MulTIMaskedN mul2 (
    .io_x_0     (e_0[3:0]           ), //i
    .io_x_1     (e_1[3:0]           ), //i
    .io_x_2     (e_2[3:0]           ), //i
    .io_x_3     (e_3[3:0]           ), //i
    .io_x_4     (e_4[3:0]           ), //i
    .io_x_5     (e_5[3:0]           ), //i
    .io_x_6     (e_6[3:0]           ), //i
    .io_x_7     (e_7[3:0]           ), //i
    .io_x_8     (e_8[3:0]           ), //i
    .io_x_9     (e_9[3:0]           ), //i
    .io_x_10    (e_10[3:0]          ), //i
    .io_x_11    (e_11[3:0]          ), //i
    .io_x_12    (e_12[3:0]          ), //i
    .io_y_0     (b_0[3:0]           ), //i
    .io_y_1     (b_1[3:0]           ), //i
    .io_y_2     (b_2[3:0]           ), //i
    .io_y_3     (b_3[3:0]           ), //i
    .io_y_4     (b_4[3:0]           ), //i
    .io_y_5     (b_5[3:0]           ), //i
    .io_y_6     (b_6[3:0]           ), //i
    .io_y_7     (b_7[3:0]           ), //i
    .io_y_8     (b_8[3:0]           ), //i
    .io_y_9     (b_9[3:0]           ), //i
    .io_y_10    (b_10[3:0]          ), //i
    .io_y_11    (b_11[3:0]          ), //i
    .io_y_12    (b_12[3:0]          ), //i
    .io_z_0     (mul2_io_z_0[3:0]   ), //o
    .io_z_1     (mul2_io_z_1[3:0]   ), //o
    .io_z_2     (mul2_io_z_2[3:0]   ), //o
    .io_z_3     (mul2_io_z_3[3:0]   ), //o
    .io_z_4     (mul2_io_z_4[3:0]   ), //o
    .io_z_5     (mul2_io_z_5[3:0]   ), //o
    .io_z_6     (mul2_io_z_6[3:0]   ), //o
    .io_z_7     (mul2_io_z_7[3:0]   ), //o
    .io_z_8     (mul2_io_z_8[3:0]   ), //o
    .io_z_9     (mul2_io_z_9[3:0]   ), //o
    .io_z_10    (mul2_io_z_10[3:0]  ), //o
    .io_z_11    (mul2_io_z_11[3:0]  ), //o
    .io_z_12    (mul2_io_z_12[3:0]  ), //o
    .clk        (clk                ), //i
    .reset      (reset              )  //i
  );
  G16MulTIMaskedN mul3 (
    .io_x_0     (e_0[3:0]           ), //i
    .io_x_1     (e_1[3:0]           ), //i
    .io_x_2     (e_2[3:0]           ), //i
    .io_x_3     (e_3[3:0]           ), //i
    .io_x_4     (e_4[3:0]           ), //i
    .io_x_5     (e_5[3:0]           ), //i
    .io_x_6     (e_6[3:0]           ), //i
    .io_x_7     (e_7[3:0]           ), //i
    .io_x_8     (e_8[3:0]           ), //i
    .io_x_9     (e_9[3:0]           ), //i
    .io_x_10    (e_10[3:0]          ), //i
    .io_x_11    (e_11[3:0]          ), //i
    .io_x_12    (e_12[3:0]          ), //i
    .io_y_0     (a_0[3:0]           ), //i
    .io_y_1     (a_1[3:0]           ), //i
    .io_y_2     (a_2[3:0]           ), //i
    .io_y_3     (a_3[3:0]           ), //i
    .io_y_4     (a_4[3:0]           ), //i
    .io_y_5     (a_5[3:0]           ), //i
    .io_y_6     (a_6[3:0]           ), //i
    .io_y_7     (a_7[3:0]           ), //i
    .io_y_8     (a_8[3:0]           ), //i
    .io_y_9     (a_9[3:0]           ), //i
    .io_y_10    (a_10[3:0]          ), //i
    .io_y_11    (a_11[3:0]          ), //i
    .io_y_12    (a_12[3:0]          ), //i
    .io_z_0     (mul3_io_z_0[3:0]   ), //o
    .io_z_1     (mul3_io_z_1[3:0]   ), //o
    .io_z_2     (mul3_io_z_2[3:0]   ), //o
    .io_z_3     (mul3_io_z_3[3:0]   ), //o
    .io_z_4     (mul3_io_z_4[3:0]   ), //o
    .io_z_5     (mul3_io_z_5[3:0]   ), //o
    .io_z_6     (mul3_io_z_6[3:0]   ), //o
    .io_z_7     (mul3_io_z_7[3:0]   ), //o
    .io_z_8     (mul3_io_z_8[3:0]   ), //o
    .io_z_9     (mul3_io_z_9[3:0]   ), //o
    .io_z_10    (mul3_io_z_10[3:0]  ), //o
    .io_z_11    (mul3_io_z_11[3:0]  ), //o
    .io_z_12    (mul3_io_z_12[3:0]  ), //o
    .clk        (clk                ), //i
    .reset      (reset              )  //i
  );
  G16InvTIMaskedN inv (
    .io_x_0     (inv_io_x_0[3:0]   ), //i
    .io_x_1     (inv_io_x_1[3:0]   ), //i
    .io_x_2     (inv_io_x_2[3:0]   ), //i
    .io_x_3     (inv_io_x_3[3:0]   ), //i
    .io_x_4     (inv_io_x_4[3:0]   ), //i
    .io_x_5     (inv_io_x_5[3:0]   ), //i
    .io_x_6     (inv_io_x_6[3:0]   ), //i
    .io_x_7     (inv_io_x_7[3:0]   ), //i
    .io_x_8     (inv_io_x_8[3:0]   ), //i
    .io_x_9     (inv_io_x_9[3:0]   ), //i
    .io_x_10    (inv_io_x_10[3:0]  ), //i
    .io_x_11    (inv_io_x_11[3:0]  ), //i
    .io_x_12    (inv_io_x_12[3:0]  ), //i
    .io_z_0     (inv_io_z_0[3:0]   ), //o
    .io_z_1     (inv_io_z_1[3:0]   ), //o
    .io_z_2     (inv_io_z_2[3:0]   ), //o
    .io_z_3     (inv_io_z_3[3:0]   ), //o
    .io_z_4     (inv_io_z_4[3:0]   ), //o
    .io_z_5     (inv_io_z_5[3:0]   ), //o
    .io_z_6     (inv_io_z_6[3:0]   ), //o
    .io_z_7     (inv_io_z_7[3:0]   ), //o
    .io_z_8     (inv_io_z_8[3:0]   ), //o
    .io_z_9     (inv_io_z_9[3:0]   ), //o
    .io_z_10    (inv_io_z_10[3:0]  ), //o
    .io_z_11    (inv_io_z_11[3:0]  ), //o
    .io_z_12    (inv_io_z_12[3:0]  ), //o
    .clk        (clk               ), //i
    .reset      (reset             )  //i
  );
  G16SqSc g16SqSc_13 (
    .io_t    (f_0[3:0]              ), //i
    .io_x    (g16SqSc_13_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_14 (
    .io_t    (f_1[3:0]              ), //i
    .io_x    (g16SqSc_14_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_15 (
    .io_t    (f_2[3:0]              ), //i
    .io_x    (g16SqSc_15_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_16 (
    .io_t    (f_3[3:0]              ), //i
    .io_x    (g16SqSc_16_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_17 (
    .io_t    (f_4[3:0]              ), //i
    .io_x    (g16SqSc_17_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_18 (
    .io_t    (f_5[3:0]              ), //i
    .io_x    (g16SqSc_18_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_19 (
    .io_t    (f_6[3:0]              ), //i
    .io_x    (g16SqSc_19_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_20 (
    .io_t    (f_7[3:0]              ), //i
    .io_x    (g16SqSc_20_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_21 (
    .io_t    (f_8[3:0]              ), //i
    .io_x    (g16SqSc_21_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_22 (
    .io_t    (f_9[3:0]              ), //i
    .io_x    (g16SqSc_22_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_23 (
    .io_t    (f_10[3:0]             ), //i
    .io_x    (g16SqSc_23_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_24 (
    .io_t    (f_11[3:0]             ), //i
    .io_x    (g16SqSc_24_io_x[3:0]  )  //o
  );
  G16SqSc g16SqSc_25 (
    .io_t    (f_12[3:0]             ), //i
    .io_x    (g16SqSc_25_io_x[3:0]  )  //o
  );
  assign dummy = 1'b0;
  assign a_0 = io_x_0[7 : 4];
  assign b_0 = io_x_0[3 : 0];
  assign a_1 = io_x_1[7 : 4];
  assign b_1 = io_x_1[3 : 0];
  assign a_2 = io_x_2[7 : 4];
  assign b_2 = io_x_2[3 : 0];
  assign a_3 = io_x_3[7 : 4];
  assign b_3 = io_x_3[3 : 0];
  assign a_4 = io_x_4[7 : 4];
  assign b_4 = io_x_4[3 : 0];
  assign a_5 = io_x_5[7 : 4];
  assign b_5 = io_x_5[3 : 0];
  assign a_6 = io_x_6[7 : 4];
  assign b_6 = io_x_6[3 : 0];
  assign a_7 = io_x_7[7 : 4];
  assign b_7 = io_x_7[3 : 0];
  assign a_8 = io_x_8[7 : 4];
  assign b_8 = io_x_8[3 : 0];
  assign a_9 = io_x_9[7 : 4];
  assign b_9 = io_x_9[3 : 0];
  assign a_10 = io_x_10[7 : 4];
  assign b_10 = io_x_10[3 : 0];
  assign a_11 = io_x_11[7 : 4];
  assign b_11 = io_x_11[3 : 0];
  assign a_12 = io_x_12[7 : 4];
  assign b_12 = io_x_12[3 : 0];
  assign f_0 = (a_0 ^ b_0);
  assign f_1 = (a_1 ^ b_1);
  assign f_2 = (a_2 ^ b_2);
  assign f_3 = (a_3 ^ b_3);
  assign f_4 = (a_4 ^ b_4);
  assign f_5 = (a_5 ^ b_5);
  assign f_6 = (a_6 ^ b_6);
  assign f_7 = (a_7 ^ b_7);
  assign f_8 = (a_8 ^ b_8);
  assign f_9 = (a_9 ^ b_9);
  assign f_10 = (a_10 ^ b_10);
  assign f_11 = (a_11 ^ b_11);
  assign f_12 = (a_12 ^ b_12);
  assign c_0 = g16SqSc_13_io_x;
  assign c_1 = g16SqSc_14_io_x;
  assign c_2 = g16SqSc_15_io_x;
  assign c_3 = g16SqSc_16_io_x;
  assign c_4 = g16SqSc_17_io_x;
  assign c_5 = g16SqSc_18_io_x;
  assign c_6 = g16SqSc_19_io_x;
  assign c_7 = g16SqSc_20_io_x;
  assign c_8 = g16SqSc_21_io_x;
  assign c_9 = g16SqSc_22_io_x;
  assign c_10 = g16SqSc_23_io_x;
  assign c_11 = g16SqSc_24_io_x;
  assign c_12 = g16SqSc_25_io_x;
  assign d_0 = mul1_io_z_0;
  assign d_1 = mul1_io_z_1;
  assign d_2 = mul1_io_z_2;
  assign d_3 = mul1_io_z_3;
  assign d_4 = mul1_io_z_4;
  assign d_5 = mul1_io_z_5;
  assign d_6 = mul1_io_z_6;
  assign d_7 = mul1_io_z_7;
  assign d_8 = mul1_io_z_8;
  assign d_9 = mul1_io_z_9;
  assign d_10 = mul1_io_z_10;
  assign d_11 = mul1_io_z_11;
  assign d_12 = mul1_io_z_12;
  assign inv_io_x_0 = (c_0 ^ d_0);
  assign inv_io_x_1 = (c_1 ^ d_1);
  assign inv_io_x_2 = (c_2 ^ d_2);
  assign inv_io_x_3 = (c_3 ^ d_3);
  assign inv_io_x_4 = (c_4 ^ d_4);
  assign inv_io_x_5 = (c_5 ^ d_5);
  assign inv_io_x_6 = (c_6 ^ d_6);
  assign inv_io_x_7 = (c_7 ^ d_7);
  assign inv_io_x_8 = (c_8 ^ d_8);
  assign inv_io_x_9 = (c_9 ^ d_9);
  assign inv_io_x_10 = (c_10 ^ d_10);
  assign inv_io_x_11 = (c_11 ^ d_11);
  assign inv_io_x_12 = (c_12 ^ d_12);
  assign e_0 = inv_io_z_0;
  assign e_1 = inv_io_z_1;
  assign e_2 = inv_io_z_2;
  assign e_3 = inv_io_z_3;
  assign e_4 = inv_io_z_4;
  assign e_5 = inv_io_z_5;
  assign e_6 = inv_io_z_6;
  assign e_7 = inv_io_z_7;
  assign e_8 = inv_io_z_8;
  assign e_9 = inv_io_z_9;
  assign e_10 = inv_io_z_10;
  assign e_11 = inv_io_z_11;
  assign e_12 = inv_io_z_12;
  assign p_0 = mul2_io_z_0;
  assign p_1 = mul2_io_z_1;
  assign p_2 = mul2_io_z_2;
  assign p_3 = mul2_io_z_3;
  assign p_4 = mul2_io_z_4;
  assign p_5 = mul2_io_z_5;
  assign p_6 = mul2_io_z_6;
  assign p_7 = mul2_io_z_7;
  assign p_8 = mul2_io_z_8;
  assign p_9 = mul2_io_z_9;
  assign p_10 = mul2_io_z_10;
  assign p_11 = mul2_io_z_11;
  assign p_12 = mul2_io_z_12;
  assign q_0 = mul3_io_z_0;
  assign q_1 = mul3_io_z_1;
  assign q_2 = mul3_io_z_2;
  assign q_3 = mul3_io_z_3;
  assign q_4 = mul3_io_z_4;
  assign q_5 = mul3_io_z_5;
  assign q_6 = mul3_io_z_6;
  assign q_7 = mul3_io_z_7;
  assign q_8 = mul3_io_z_8;
  assign q_9 = mul3_io_z_9;
  assign q_10 = mul3_io_z_10;
  assign q_11 = mul3_io_z_11;
  assign q_12 = mul3_io_z_12;
  assign io_z_0 = {p_0,q_0};
  assign io_z_1 = {p_1,q_1};
  assign io_z_2 = {p_2,q_2};
  assign io_z_3 = {p_3,q_3};
  assign io_z_4 = {p_4,q_4};
  assign io_z_5 = {p_5,q_5};
  assign io_z_6 = {p_6,q_6};
  assign io_z_7 = {p_7,q_7};
  assign io_z_8 = {p_8,q_8};
  assign io_z_9 = {p_9,q_9};
  assign io_z_10 = {p_10,q_10};
  assign io_z_11 = {p_11,q_11};
  assign io_z_12 = {p_12,q_12};

endmodule

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

//G16SqSc replaced by G16SqSc

module G16SqSc (
  input      [3:0]    io_t,
  output     [3:0]    io_x
);

  wire       [1:0]    square1_io_t;
  wire       [1:0]    square1_io_x;
  wire       [1:0]    square2_io_x;
  wire       [1:0]    scale_io_x;
  wire       [1:0]    a;
  wire       [1:0]    b;
  wire       [1:0]    c;
  wire       [1:0]    p;
  wire       [1:0]    q;

  G4Sq square1 (
    .io_t    (square1_io_t[1:0]  ), //i
    .io_x    (square1_io_x[1:0]  )  //o
  );
  G4Sq square2 (
    .io_t    (b[1:0]             ), //i
    .io_x    (square2_io_x[1:0]  )  //o
  );
  G4ScaleN2 scale (
    .io_t    (c[1:0]           ), //i
    .io_x    (scale_io_x[1:0]  )  //o
  );
  assign square1_io_t = (a ^ b);
  assign p = square1_io_x;
  assign c = square2_io_x;
  assign q = scale_io_x;
  assign a = io_t[3 : 2];
  assign b = io_t[1 : 0];
  assign io_x = {p,q};

endmodule

module G16InvTIMaskedN (
  input      [3:0]    io_x_0,
  input      [3:0]    io_x_1,
  input      [3:0]    io_x_2,
  input      [3:0]    io_x_3,
  input      [3:0]    io_x_4,
  input      [3:0]    io_x_5,
  input      [3:0]    io_x_6,
  input      [3:0]    io_x_7,
  input      [3:0]    io_x_8,
  input      [3:0]    io_x_9,
  input      [3:0]    io_x_10,
  input      [3:0]    io_x_11,
  input      [3:0]    io_x_12,
  output     [3:0]    io_z_0,
  output     [3:0]    io_z_1,
  output     [3:0]    io_z_2,
  output     [3:0]    io_z_3,
  output     [3:0]    io_z_4,
  output     [3:0]    io_z_5,
  output     [3:0]    io_z_6,
  output     [3:0]    io_z_7,
  output     [3:0]    io_z_8,
  output     [3:0]    io_z_9,
  output     [3:0]    io_z_10,
  output     [3:0]    io_z_11,
  output     [3:0]    io_z_12,
  input               clk,
  input               reset
);

  wire       [1:0]    g4Sq_65_io_t;
  wire       [1:0]    g4Sq_66_io_t;
  wire       [1:0]    g4Sq_67_io_t;
  wire       [1:0]    g4Sq_68_io_t;
  wire       [1:0]    g4Sq_69_io_t;
  wire       [1:0]    g4Sq_70_io_t;
  wire       [1:0]    g4Sq_71_io_t;
  wire       [1:0]    g4Sq_72_io_t;
  wire       [1:0]    g4Sq_73_io_t;
  wire       [1:0]    g4Sq_74_io_t;
  wire       [1:0]    g4Sq_75_io_t;
  wire       [1:0]    g4Sq_76_io_t;
  wire       [1:0]    g4Sq_77_io_t;
  wire       [1:0]    mul1_io_z_0;
  wire       [1:0]    mul1_io_z_1;
  wire       [1:0]    mul1_io_z_2;
  wire       [1:0]    mul1_io_z_3;
  wire       [1:0]    mul1_io_z_4;
  wire       [1:0]    mul1_io_z_5;
  wire       [1:0]    mul1_io_z_6;
  wire       [1:0]    mul1_io_z_7;
  wire       [1:0]    mul1_io_z_8;
  wire       [1:0]    mul1_io_z_9;
  wire       [1:0]    mul1_io_z_10;
  wire       [1:0]    mul1_io_z_11;
  wire       [1:0]    mul1_io_z_12;
  wire       [1:0]    mul2_io_z_0;
  wire       [1:0]    mul2_io_z_1;
  wire       [1:0]    mul2_io_z_2;
  wire       [1:0]    mul2_io_z_3;
  wire       [1:0]    mul2_io_z_4;
  wire       [1:0]    mul2_io_z_5;
  wire       [1:0]    mul2_io_z_6;
  wire       [1:0]    mul2_io_z_7;
  wire       [1:0]    mul2_io_z_8;
  wire       [1:0]    mul2_io_z_9;
  wire       [1:0]    mul2_io_z_10;
  wire       [1:0]    mul2_io_z_11;
  wire       [1:0]    mul2_io_z_12;
  wire       [1:0]    mul3_io_z_0;
  wire       [1:0]    mul3_io_z_1;
  wire       [1:0]    mul3_io_z_2;
  wire       [1:0]    mul3_io_z_3;
  wire       [1:0]    mul3_io_z_4;
  wire       [1:0]    mul3_io_z_5;
  wire       [1:0]    mul3_io_z_6;
  wire       [1:0]    mul3_io_z_7;
  wire       [1:0]    mul3_io_z_8;
  wire       [1:0]    mul3_io_z_9;
  wire       [1:0]    mul3_io_z_10;
  wire       [1:0]    mul3_io_z_11;
  wire       [1:0]    mul3_io_z_12;
  wire       [1:0]    g4Sq_52_io_x;
  wire       [1:0]    g4ScaleN_52_io_x;
  wire       [1:0]    g4Sq_53_io_x;
  wire       [1:0]    g4ScaleN_53_io_x;
  wire       [1:0]    g4Sq_54_io_x;
  wire       [1:0]    g4ScaleN_54_io_x;
  wire       [1:0]    g4Sq_55_io_x;
  wire       [1:0]    g4ScaleN_55_io_x;
  wire       [1:0]    g4Sq_56_io_x;
  wire       [1:0]    g4ScaleN_56_io_x;
  wire       [1:0]    g4Sq_57_io_x;
  wire       [1:0]    g4ScaleN_57_io_x;
  wire       [1:0]    g4Sq_58_io_x;
  wire       [1:0]    g4ScaleN_58_io_x;
  wire       [1:0]    g4Sq_59_io_x;
  wire       [1:0]    g4ScaleN_59_io_x;
  wire       [1:0]    g4Sq_60_io_x;
  wire       [1:0]    g4ScaleN_60_io_x;
  wire       [1:0]    g4Sq_61_io_x;
  wire       [1:0]    g4ScaleN_61_io_x;
  wire       [1:0]    g4Sq_62_io_x;
  wire       [1:0]    g4ScaleN_62_io_x;
  wire       [1:0]    g4Sq_63_io_x;
  wire       [1:0]    g4ScaleN_63_io_x;
  wire       [1:0]    g4Sq_64_io_x;
  wire       [1:0]    g4ScaleN_64_io_x;
  wire       [1:0]    g4Sq_65_io_x;
  wire       [1:0]    g4Sq_66_io_x;
  wire       [1:0]    g4Sq_67_io_x;
  wire       [1:0]    g4Sq_68_io_x;
  wire       [1:0]    g4Sq_69_io_x;
  wire       [1:0]    g4Sq_70_io_x;
  wire       [1:0]    g4Sq_71_io_x;
  wire       [1:0]    g4Sq_72_io_x;
  wire       [1:0]    g4Sq_73_io_x;
  wire       [1:0]    g4Sq_74_io_x;
  wire       [1:0]    g4Sq_75_io_x;
  wire       [1:0]    g4Sq_76_io_x;
  wire       [1:0]    g4Sq_77_io_x;
  wire                dummy;
  wire       [1:0]    a_0;
  wire       [1:0]    a_1;
  wire       [1:0]    a_2;
  wire       [1:0]    a_3;
  wire       [1:0]    a_4;
  wire       [1:0]    a_5;
  wire       [1:0]    a_6;
  wire       [1:0]    a_7;
  wire       [1:0]    a_8;
  wire       [1:0]    a_9;
  wire       [1:0]    a_10;
  wire       [1:0]    a_11;
  wire       [1:0]    a_12;
  wire       [1:0]    b_0;
  wire       [1:0]    b_1;
  wire       [1:0]    b_2;
  wire       [1:0]    b_3;
  wire       [1:0]    b_4;
  wire       [1:0]    b_5;
  wire       [1:0]    b_6;
  wire       [1:0]    b_7;
  wire       [1:0]    b_8;
  wire       [1:0]    b_9;
  wire       [1:0]    b_10;
  wire       [1:0]    b_11;
  wire       [1:0]    b_12;
  wire       [1:0]    c_0;
  wire       [1:0]    c_1;
  wire       [1:0]    c_2;
  wire       [1:0]    c_3;
  wire       [1:0]    c_4;
  wire       [1:0]    c_5;
  wire       [1:0]    c_6;
  wire       [1:0]    c_7;
  wire       [1:0]    c_8;
  wire       [1:0]    c_9;
  wire       [1:0]    c_10;
  wire       [1:0]    c_11;
  wire       [1:0]    c_12;
  wire       [1:0]    d_0;
  wire       [1:0]    d_1;
  wire       [1:0]    d_2;
  wire       [1:0]    d_3;
  wire       [1:0]    d_4;
  wire       [1:0]    d_5;
  wire       [1:0]    d_6;
  wire       [1:0]    d_7;
  wire       [1:0]    d_8;
  wire       [1:0]    d_9;
  wire       [1:0]    d_10;
  wire       [1:0]    d_11;
  wire       [1:0]    d_12;
  wire       [1:0]    e_0;
  wire       [1:0]    e_1;
  wire       [1:0]    e_2;
  wire       [1:0]    e_3;
  wire       [1:0]    e_4;
  wire       [1:0]    e_5;
  wire       [1:0]    e_6;
  wire       [1:0]    e_7;
  wire       [1:0]    e_8;
  wire       [1:0]    e_9;
  wire       [1:0]    e_10;
  wire       [1:0]    e_11;
  wire       [1:0]    e_12;
  wire       [1:0]    f_0;
  wire       [1:0]    f_1;
  wire       [1:0]    f_2;
  wire       [1:0]    f_3;
  wire       [1:0]    f_4;
  wire       [1:0]    f_5;
  wire       [1:0]    f_6;
  wire       [1:0]    f_7;
  wire       [1:0]    f_8;
  wire       [1:0]    f_9;
  wire       [1:0]    f_10;
  wire       [1:0]    f_11;
  wire       [1:0]    f_12;
  wire       [1:0]    p_0;
  wire       [1:0]    p_1;
  wire       [1:0]    p_2;
  wire       [1:0]    p_3;
  wire       [1:0]    p_4;
  wire       [1:0]    p_5;
  wire       [1:0]    p_6;
  wire       [1:0]    p_7;
  wire       [1:0]    p_8;
  wire       [1:0]    p_9;
  wire       [1:0]    p_10;
  wire       [1:0]    p_11;
  wire       [1:0]    p_12;
  wire       [1:0]    q_0;
  wire       [1:0]    q_1;
  wire       [1:0]    q_2;
  wire       [1:0]    q_3;
  wire       [1:0]    q_4;
  wire       [1:0]    q_5;
  wire       [1:0]    q_6;
  wire       [1:0]    q_7;
  wire       [1:0]    q_8;
  wire       [1:0]    q_9;
  wire       [1:0]    q_10;
  wire       [1:0]    q_11;
  wire       [1:0]    q_12;

  G4MulTIMaskedN mul1 (
    .io_x_0     (a_0[1:0]           ), //i
    .io_x_1     (a_1[1:0]           ), //i
    .io_x_2     (a_2[1:0]           ), //i
    .io_x_3     (a_3[1:0]           ), //i
    .io_x_4     (a_4[1:0]           ), //i
    .io_x_5     (a_5[1:0]           ), //i
    .io_x_6     (a_6[1:0]           ), //i
    .io_x_7     (a_7[1:0]           ), //i
    .io_x_8     (a_8[1:0]           ), //i
    .io_x_9     (a_9[1:0]           ), //i
    .io_x_10    (a_10[1:0]          ), //i
    .io_x_11    (a_11[1:0]          ), //i
    .io_x_12    (a_12[1:0]          ), //i
    .io_y_0     (b_0[1:0]           ), //i
    .io_y_1     (b_1[1:0]           ), //i
    .io_y_2     (b_2[1:0]           ), //i
    .io_y_3     (b_3[1:0]           ), //i
    .io_y_4     (b_4[1:0]           ), //i
    .io_y_5     (b_5[1:0]           ), //i
    .io_y_6     (b_6[1:0]           ), //i
    .io_y_7     (b_7[1:0]           ), //i
    .io_y_8     (b_8[1:0]           ), //i
    .io_y_9     (b_9[1:0]           ), //i
    .io_y_10    (b_10[1:0]          ), //i
    .io_y_11    (b_11[1:0]          ), //i
    .io_y_12    (b_12[1:0]          ), //i
    .io_z_0     (mul1_io_z_0[1:0]   ), //o
    .io_z_1     (mul1_io_z_1[1:0]   ), //o
    .io_z_2     (mul1_io_z_2[1:0]   ), //o
    .io_z_3     (mul1_io_z_3[1:0]   ), //o
    .io_z_4     (mul1_io_z_4[1:0]   ), //o
    .io_z_5     (mul1_io_z_5[1:0]   ), //o
    .io_z_6     (mul1_io_z_6[1:0]   ), //o
    .io_z_7     (mul1_io_z_7[1:0]   ), //o
    .io_z_8     (mul1_io_z_8[1:0]   ), //o
    .io_z_9     (mul1_io_z_9[1:0]   ), //o
    .io_z_10    (mul1_io_z_10[1:0]  ), //o
    .io_z_11    (mul1_io_z_11[1:0]  ), //o
    .io_z_12    (mul1_io_z_12[1:0]  ), //o
    .clk        (clk                ), //i
    .reset      (reset              )  //i
  );
  G4MulTIMaskedN mul2 (
    .io_x_0     (e_0[1:0]           ), //i
    .io_x_1     (e_1[1:0]           ), //i
    .io_x_2     (e_2[1:0]           ), //i
    .io_x_3     (e_3[1:0]           ), //i
    .io_x_4     (e_4[1:0]           ), //i
    .io_x_5     (e_5[1:0]           ), //i
    .io_x_6     (e_6[1:0]           ), //i
    .io_x_7     (e_7[1:0]           ), //i
    .io_x_8     (e_8[1:0]           ), //i
    .io_x_9     (e_9[1:0]           ), //i
    .io_x_10    (e_10[1:0]          ), //i
    .io_x_11    (e_11[1:0]          ), //i
    .io_x_12    (e_12[1:0]          ), //i
    .io_y_0     (b_0[1:0]           ), //i
    .io_y_1     (b_1[1:0]           ), //i
    .io_y_2     (b_2[1:0]           ), //i
    .io_y_3     (b_3[1:0]           ), //i
    .io_y_4     (b_4[1:0]           ), //i
    .io_y_5     (b_5[1:0]           ), //i
    .io_y_6     (b_6[1:0]           ), //i
    .io_y_7     (b_7[1:0]           ), //i
    .io_y_8     (b_8[1:0]           ), //i
    .io_y_9     (b_9[1:0]           ), //i
    .io_y_10    (b_10[1:0]          ), //i
    .io_y_11    (b_11[1:0]          ), //i
    .io_y_12    (b_12[1:0]          ), //i
    .io_z_0     (mul2_io_z_0[1:0]   ), //o
    .io_z_1     (mul2_io_z_1[1:0]   ), //o
    .io_z_2     (mul2_io_z_2[1:0]   ), //o
    .io_z_3     (mul2_io_z_3[1:0]   ), //o
    .io_z_4     (mul2_io_z_4[1:0]   ), //o
    .io_z_5     (mul2_io_z_5[1:0]   ), //o
    .io_z_6     (mul2_io_z_6[1:0]   ), //o
    .io_z_7     (mul2_io_z_7[1:0]   ), //o
    .io_z_8     (mul2_io_z_8[1:0]   ), //o
    .io_z_9     (mul2_io_z_9[1:0]   ), //o
    .io_z_10    (mul2_io_z_10[1:0]  ), //o
    .io_z_11    (mul2_io_z_11[1:0]  ), //o
    .io_z_12    (mul2_io_z_12[1:0]  ), //o
    .clk        (clk                ), //i
    .reset      (reset              )  //i
  );
  G4MulTIMaskedN mul3 (
    .io_x_0     (e_0[1:0]           ), //i
    .io_x_1     (e_1[1:0]           ), //i
    .io_x_2     (e_2[1:0]           ), //i
    .io_x_3     (e_3[1:0]           ), //i
    .io_x_4     (e_4[1:0]           ), //i
    .io_x_5     (e_5[1:0]           ), //i
    .io_x_6     (e_6[1:0]           ), //i
    .io_x_7     (e_7[1:0]           ), //i
    .io_x_8     (e_8[1:0]           ), //i
    .io_x_9     (e_9[1:0]           ), //i
    .io_x_10    (e_10[1:0]          ), //i
    .io_x_11    (e_11[1:0]          ), //i
    .io_x_12    (e_12[1:0]          ), //i
    .io_y_0     (a_0[1:0]           ), //i
    .io_y_1     (a_1[1:0]           ), //i
    .io_y_2     (a_2[1:0]           ), //i
    .io_y_3     (a_3[1:0]           ), //i
    .io_y_4     (a_4[1:0]           ), //i
    .io_y_5     (a_5[1:0]           ), //i
    .io_y_6     (a_6[1:0]           ), //i
    .io_y_7     (a_7[1:0]           ), //i
    .io_y_8     (a_8[1:0]           ), //i
    .io_y_9     (a_9[1:0]           ), //i
    .io_y_10    (a_10[1:0]          ), //i
    .io_y_11    (a_11[1:0]          ), //i
    .io_y_12    (a_12[1:0]          ), //i
    .io_z_0     (mul3_io_z_0[1:0]   ), //o
    .io_z_1     (mul3_io_z_1[1:0]   ), //o
    .io_z_2     (mul3_io_z_2[1:0]   ), //o
    .io_z_3     (mul3_io_z_3[1:0]   ), //o
    .io_z_4     (mul3_io_z_4[1:0]   ), //o
    .io_z_5     (mul3_io_z_5[1:0]   ), //o
    .io_z_6     (mul3_io_z_6[1:0]   ), //o
    .io_z_7     (mul3_io_z_7[1:0]   ), //o
    .io_z_8     (mul3_io_z_8[1:0]   ), //o
    .io_z_9     (mul3_io_z_9[1:0]   ), //o
    .io_z_10    (mul3_io_z_10[1:0]  ), //o
    .io_z_11    (mul3_io_z_11[1:0]  ), //o
    .io_z_12    (mul3_io_z_12[1:0]  ), //o
    .clk        (clk                ), //i
    .reset      (reset              )  //i
  );
  G4Sq g4Sq_52 (
    .io_t    (f_0[1:0]           ), //i
    .io_x    (g4Sq_52_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_52 (
    .io_t    (g4Sq_52_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_52_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_53 (
    .io_t    (f_1[1:0]           ), //i
    .io_x    (g4Sq_53_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_53 (
    .io_t    (g4Sq_53_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_53_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_54 (
    .io_t    (f_2[1:0]           ), //i
    .io_x    (g4Sq_54_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_54 (
    .io_t    (g4Sq_54_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_54_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_55 (
    .io_t    (f_3[1:0]           ), //i
    .io_x    (g4Sq_55_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_55 (
    .io_t    (g4Sq_55_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_55_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_56 (
    .io_t    (f_4[1:0]           ), //i
    .io_x    (g4Sq_56_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_56 (
    .io_t    (g4Sq_56_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_56_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_57 (
    .io_t    (f_5[1:0]           ), //i
    .io_x    (g4Sq_57_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_57 (
    .io_t    (g4Sq_57_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_57_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_58 (
    .io_t    (f_6[1:0]           ), //i
    .io_x    (g4Sq_58_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_58 (
    .io_t    (g4Sq_58_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_58_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_59 (
    .io_t    (f_7[1:0]           ), //i
    .io_x    (g4Sq_59_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_59 (
    .io_t    (g4Sq_59_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_59_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_60 (
    .io_t    (f_8[1:0]           ), //i
    .io_x    (g4Sq_60_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_60 (
    .io_t    (g4Sq_60_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_60_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_61 (
    .io_t    (f_9[1:0]           ), //i
    .io_x    (g4Sq_61_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_61 (
    .io_t    (g4Sq_61_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_61_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_62 (
    .io_t    (f_10[1:0]          ), //i
    .io_x    (g4Sq_62_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_62 (
    .io_t    (g4Sq_62_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_62_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_63 (
    .io_t    (f_11[1:0]          ), //i
    .io_x    (g4Sq_63_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_63 (
    .io_t    (g4Sq_63_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_63_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_64 (
    .io_t    (f_12[1:0]          ), //i
    .io_x    (g4Sq_64_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_64 (
    .io_t    (g4Sq_64_io_x[1:0]      ), //i
    .io_x    (g4ScaleN_64_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_65 (
    .io_t    (g4Sq_65_io_t[1:0]  ), //i
    .io_x    (g4Sq_65_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_66 (
    .io_t    (g4Sq_66_io_t[1:0]  ), //i
    .io_x    (g4Sq_66_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_67 (
    .io_t    (g4Sq_67_io_t[1:0]  ), //i
    .io_x    (g4Sq_67_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_68 (
    .io_t    (g4Sq_68_io_t[1:0]  ), //i
    .io_x    (g4Sq_68_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_69 (
    .io_t    (g4Sq_69_io_t[1:0]  ), //i
    .io_x    (g4Sq_69_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_70 (
    .io_t    (g4Sq_70_io_t[1:0]  ), //i
    .io_x    (g4Sq_70_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_71 (
    .io_t    (g4Sq_71_io_t[1:0]  ), //i
    .io_x    (g4Sq_71_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_72 (
    .io_t    (g4Sq_72_io_t[1:0]  ), //i
    .io_x    (g4Sq_72_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_73 (
    .io_t    (g4Sq_73_io_t[1:0]  ), //i
    .io_x    (g4Sq_73_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_74 (
    .io_t    (g4Sq_74_io_t[1:0]  ), //i
    .io_x    (g4Sq_74_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_75 (
    .io_t    (g4Sq_75_io_t[1:0]  ), //i
    .io_x    (g4Sq_75_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_76 (
    .io_t    (g4Sq_76_io_t[1:0]  ), //i
    .io_x    (g4Sq_76_io_x[1:0]  )  //o
  );
  G4Sq g4Sq_77 (
    .io_t    (g4Sq_77_io_t[1:0]  ), //i
    .io_x    (g4Sq_77_io_x[1:0]  )  //o
  );
  assign dummy = 1'b0;
  assign a_0 = io_x_0[3 : 2];
  assign b_0 = io_x_0[1 : 0];
  assign a_1 = io_x_1[3 : 2];
  assign b_1 = io_x_1[1 : 0];
  assign a_2 = io_x_2[3 : 2];
  assign b_2 = io_x_2[1 : 0];
  assign a_3 = io_x_3[3 : 2];
  assign b_3 = io_x_3[1 : 0];
  assign a_4 = io_x_4[3 : 2];
  assign b_4 = io_x_4[1 : 0];
  assign a_5 = io_x_5[3 : 2];
  assign b_5 = io_x_5[1 : 0];
  assign a_6 = io_x_6[3 : 2];
  assign b_6 = io_x_6[1 : 0];
  assign a_7 = io_x_7[3 : 2];
  assign b_7 = io_x_7[1 : 0];
  assign a_8 = io_x_8[3 : 2];
  assign b_8 = io_x_8[1 : 0];
  assign a_9 = io_x_9[3 : 2];
  assign b_9 = io_x_9[1 : 0];
  assign a_10 = io_x_10[3 : 2];
  assign b_10 = io_x_10[1 : 0];
  assign a_11 = io_x_11[3 : 2];
  assign b_11 = io_x_11[1 : 0];
  assign a_12 = io_x_12[3 : 2];
  assign b_12 = io_x_12[1 : 0];
  assign f_0 = (a_0 ^ b_0);
  assign f_1 = (a_1 ^ b_1);
  assign f_2 = (a_2 ^ b_2);
  assign f_3 = (a_3 ^ b_3);
  assign f_4 = (a_4 ^ b_4);
  assign f_5 = (a_5 ^ b_5);
  assign f_6 = (a_6 ^ b_6);
  assign f_7 = (a_7 ^ b_7);
  assign f_8 = (a_8 ^ b_8);
  assign f_9 = (a_9 ^ b_9);
  assign f_10 = (a_10 ^ b_10);
  assign f_11 = (a_11 ^ b_11);
  assign f_12 = (a_12 ^ b_12);
  assign d_0 = mul1_io_z_0;
  assign d_1 = mul1_io_z_1;
  assign d_2 = mul1_io_z_2;
  assign d_3 = mul1_io_z_3;
  assign d_4 = mul1_io_z_4;
  assign d_5 = mul1_io_z_5;
  assign d_6 = mul1_io_z_6;
  assign d_7 = mul1_io_z_7;
  assign d_8 = mul1_io_z_8;
  assign d_9 = mul1_io_z_9;
  assign d_10 = mul1_io_z_10;
  assign d_11 = mul1_io_z_11;
  assign d_12 = mul1_io_z_12;
  assign c_0 = g4ScaleN_52_io_x;
  assign c_1 = g4ScaleN_53_io_x;
  assign c_2 = g4ScaleN_54_io_x;
  assign c_3 = g4ScaleN_55_io_x;
  assign c_4 = g4ScaleN_56_io_x;
  assign c_5 = g4ScaleN_57_io_x;
  assign c_6 = g4ScaleN_58_io_x;
  assign c_7 = g4ScaleN_59_io_x;
  assign c_8 = g4ScaleN_60_io_x;
  assign c_9 = g4ScaleN_61_io_x;
  assign c_10 = g4ScaleN_62_io_x;
  assign c_11 = g4ScaleN_63_io_x;
  assign c_12 = g4ScaleN_64_io_x;
  assign g4Sq_65_io_t = (c_0 ^ d_0);
  assign e_0 = g4Sq_65_io_x;
  assign g4Sq_66_io_t = (c_1 ^ d_1);
  assign e_1 = g4Sq_66_io_x;
  assign g4Sq_67_io_t = (c_2 ^ d_2);
  assign e_2 = g4Sq_67_io_x;
  assign g4Sq_68_io_t = (c_3 ^ d_3);
  assign e_3 = g4Sq_68_io_x;
  assign g4Sq_69_io_t = (c_4 ^ d_4);
  assign e_4 = g4Sq_69_io_x;
  assign g4Sq_70_io_t = (c_5 ^ d_5);
  assign e_5 = g4Sq_70_io_x;
  assign g4Sq_71_io_t = (c_6 ^ d_6);
  assign e_6 = g4Sq_71_io_x;
  assign g4Sq_72_io_t = (c_7 ^ d_7);
  assign e_7 = g4Sq_72_io_x;
  assign g4Sq_73_io_t = (c_8 ^ d_8);
  assign e_8 = g4Sq_73_io_x;
  assign g4Sq_74_io_t = (c_9 ^ d_9);
  assign e_9 = g4Sq_74_io_x;
  assign g4Sq_75_io_t = (c_10 ^ d_10);
  assign e_10 = g4Sq_75_io_x;
  assign g4Sq_76_io_t = (c_11 ^ d_11);
  assign e_11 = g4Sq_76_io_x;
  assign g4Sq_77_io_t = (c_12 ^ d_12);
  assign e_12 = g4Sq_77_io_x;
  assign p_0 = mul2_io_z_0;
  assign p_1 = mul2_io_z_1;
  assign p_2 = mul2_io_z_2;
  assign p_3 = mul2_io_z_3;
  assign p_4 = mul2_io_z_4;
  assign p_5 = mul2_io_z_5;
  assign p_6 = mul2_io_z_6;
  assign p_7 = mul2_io_z_7;
  assign p_8 = mul2_io_z_8;
  assign p_9 = mul2_io_z_9;
  assign p_10 = mul2_io_z_10;
  assign p_11 = mul2_io_z_11;
  assign p_12 = mul2_io_z_12;
  assign q_0 = mul3_io_z_0;
  assign q_1 = mul3_io_z_1;
  assign q_2 = mul3_io_z_2;
  assign q_3 = mul3_io_z_3;
  assign q_4 = mul3_io_z_4;
  assign q_5 = mul3_io_z_5;
  assign q_6 = mul3_io_z_6;
  assign q_7 = mul3_io_z_7;
  assign q_8 = mul3_io_z_8;
  assign q_9 = mul3_io_z_9;
  assign q_10 = mul3_io_z_10;
  assign q_11 = mul3_io_z_11;
  assign q_12 = mul3_io_z_12;
  assign io_z_0 = {p_0,q_0};
  assign io_z_1 = {p_1,q_1};
  assign io_z_2 = {p_2,q_2};
  assign io_z_3 = {p_3,q_3};
  assign io_z_4 = {p_4,q_4};
  assign io_z_5 = {p_5,q_5};
  assign io_z_6 = {p_6,q_6};
  assign io_z_7 = {p_7,q_7};
  assign io_z_8 = {p_8,q_8};
  assign io_z_9 = {p_9,q_9};
  assign io_z_10 = {p_10,q_10};
  assign io_z_11 = {p_11,q_11};
  assign io_z_12 = {p_12,q_12};

endmodule

//G16MulTIMaskedN replaced by G16MulTIMaskedN

//G16MulTIMaskedN replaced by G16MulTIMaskedN

module G16MulTIMaskedN (
  input      [3:0]    io_x_0,
  input      [3:0]    io_x_1,
  input      [3:0]    io_x_2,
  input      [3:0]    io_x_3,
  input      [3:0]    io_x_4,
  input      [3:0]    io_x_5,
  input      [3:0]    io_x_6,
  input      [3:0]    io_x_7,
  input      [3:0]    io_x_8,
  input      [3:0]    io_x_9,
  input      [3:0]    io_x_10,
  input      [3:0]    io_x_11,
  input      [3:0]    io_x_12,
  input      [3:0]    io_y_0,
  input      [3:0]    io_y_1,
  input      [3:0]    io_y_2,
  input      [3:0]    io_y_3,
  input      [3:0]    io_y_4,
  input      [3:0]    io_y_5,
  input      [3:0]    io_y_6,
  input      [3:0]    io_y_7,
  input      [3:0]    io_y_8,
  input      [3:0]    io_y_9,
  input      [3:0]    io_y_10,
  input      [3:0]    io_y_11,
  input      [3:0]    io_y_12,
  output     [3:0]    io_z_0,
  output     [3:0]    io_z_1,
  output     [3:0]    io_z_2,
  output     [3:0]    io_z_3,
  output     [3:0]    io_z_4,
  output     [3:0]    io_z_5,
  output     [3:0]    io_z_6,
  output     [3:0]    io_z_7,
  output     [3:0]    io_z_8,
  output     [3:0]    io_z_9,
  output     [3:0]    io_z_10,
  output     [3:0]    io_z_11,
  output     [3:0]    io_z_12,
  input               clk,
  input               reset
);

  wire       [1:0]    mul1_io_x_0;
  wire       [1:0]    mul1_io_x_1;
  wire       [1:0]    mul1_io_x_2;
  wire       [1:0]    mul1_io_x_3;
  wire       [1:0]    mul1_io_x_4;
  wire       [1:0]    mul1_io_x_5;
  wire       [1:0]    mul1_io_x_6;
  wire       [1:0]    mul1_io_x_7;
  wire       [1:0]    mul1_io_x_8;
  wire       [1:0]    mul1_io_x_9;
  wire       [1:0]    mul1_io_x_10;
  wire       [1:0]    mul1_io_x_11;
  wire       [1:0]    mul1_io_x_12;
  wire       [1:0]    mul1_io_y_0;
  wire       [1:0]    mul1_io_y_1;
  wire       [1:0]    mul1_io_y_2;
  wire       [1:0]    mul1_io_y_3;
  wire       [1:0]    mul1_io_y_4;
  wire       [1:0]    mul1_io_y_5;
  wire       [1:0]    mul1_io_y_6;
  wire       [1:0]    mul1_io_y_7;
  wire       [1:0]    mul1_io_y_8;
  wire       [1:0]    mul1_io_y_9;
  wire       [1:0]    mul1_io_y_10;
  wire       [1:0]    mul1_io_y_11;
  wire       [1:0]    mul1_io_y_12;
  wire       [1:0]    mul1_io_z_0;
  wire       [1:0]    mul1_io_z_1;
  wire       [1:0]    mul1_io_z_2;
  wire       [1:0]    mul1_io_z_3;
  wire       [1:0]    mul1_io_z_4;
  wire       [1:0]    mul1_io_z_5;
  wire       [1:0]    mul1_io_z_6;
  wire       [1:0]    mul1_io_z_7;
  wire       [1:0]    mul1_io_z_8;
  wire       [1:0]    mul1_io_z_9;
  wire       [1:0]    mul1_io_z_10;
  wire       [1:0]    mul1_io_z_11;
  wire       [1:0]    mul1_io_z_12;
  wire       [1:0]    mul2_io_z_0;
  wire       [1:0]    mul2_io_z_1;
  wire       [1:0]    mul2_io_z_2;
  wire       [1:0]    mul2_io_z_3;
  wire       [1:0]    mul2_io_z_4;
  wire       [1:0]    mul2_io_z_5;
  wire       [1:0]    mul2_io_z_6;
  wire       [1:0]    mul2_io_z_7;
  wire       [1:0]    mul2_io_z_8;
  wire       [1:0]    mul2_io_z_9;
  wire       [1:0]    mul2_io_z_10;
  wire       [1:0]    mul2_io_z_11;
  wire       [1:0]    mul2_io_z_12;
  wire       [1:0]    mul3_io_z_0;
  wire       [1:0]    mul3_io_z_1;
  wire       [1:0]    mul3_io_z_2;
  wire       [1:0]    mul3_io_z_3;
  wire       [1:0]    mul3_io_z_4;
  wire       [1:0]    mul3_io_z_5;
  wire       [1:0]    mul3_io_z_6;
  wire       [1:0]    mul3_io_z_7;
  wire       [1:0]    mul3_io_z_8;
  wire       [1:0]    mul3_io_z_9;
  wire       [1:0]    mul3_io_z_10;
  wire       [1:0]    mul3_io_z_11;
  wire       [1:0]    mul3_io_z_12;
  wire       [1:0]    g4ScaleN_52_io_x;
  wire       [1:0]    g4ScaleN_53_io_x;
  wire       [1:0]    g4ScaleN_54_io_x;
  wire       [1:0]    g4ScaleN_55_io_x;
  wire       [1:0]    g4ScaleN_56_io_x;
  wire       [1:0]    g4ScaleN_57_io_x;
  wire       [1:0]    g4ScaleN_58_io_x;
  wire       [1:0]    g4ScaleN_59_io_x;
  wire       [1:0]    g4ScaleN_60_io_x;
  wire       [1:0]    g4ScaleN_61_io_x;
  wire       [1:0]    g4ScaleN_62_io_x;
  wire       [1:0]    g4ScaleN_63_io_x;
  wire       [1:0]    g4ScaleN_64_io_x;
  wire                dummy;
  wire       [1:0]    a_0;
  wire       [1:0]    a_1;
  wire       [1:0]    a_2;
  wire       [1:0]    a_3;
  wire       [1:0]    a_4;
  wire       [1:0]    a_5;
  wire       [1:0]    a_6;
  wire       [1:0]    a_7;
  wire       [1:0]    a_8;
  wire       [1:0]    a_9;
  wire       [1:0]    a_10;
  wire       [1:0]    a_11;
  wire       [1:0]    a_12;
  wire       [1:0]    b_0;
  wire       [1:0]    b_1;
  wire       [1:0]    b_2;
  wire       [1:0]    b_3;
  wire       [1:0]    b_4;
  wire       [1:0]    b_5;
  wire       [1:0]    b_6;
  wire       [1:0]    b_7;
  wire       [1:0]    b_8;
  wire       [1:0]    b_9;
  wire       [1:0]    b_10;
  wire       [1:0]    b_11;
  wire       [1:0]    b_12;
  wire       [1:0]    c_0;
  wire       [1:0]    c_1;
  wire       [1:0]    c_2;
  wire       [1:0]    c_3;
  wire       [1:0]    c_4;
  wire       [1:0]    c_5;
  wire       [1:0]    c_6;
  wire       [1:0]    c_7;
  wire       [1:0]    c_8;
  wire       [1:0]    c_9;
  wire       [1:0]    c_10;
  wire       [1:0]    c_11;
  wire       [1:0]    c_12;
  wire       [1:0]    d_0;
  wire       [1:0]    d_1;
  wire       [1:0]    d_2;
  wire       [1:0]    d_3;
  wire       [1:0]    d_4;
  wire       [1:0]    d_5;
  wire       [1:0]    d_6;
  wire       [1:0]    d_7;
  wire       [1:0]    d_8;
  wire       [1:0]    d_9;
  wire       [1:0]    d_10;
  wire       [1:0]    d_11;
  wire       [1:0]    d_12;
  wire       [1:0]    e_0;
  wire       [1:0]    e_1;
  wire       [1:0]    e_2;
  wire       [1:0]    e_3;
  wire       [1:0]    e_4;
  wire       [1:0]    e_5;
  wire       [1:0]    e_6;
  wire       [1:0]    e_7;
  wire       [1:0]    e_8;
  wire       [1:0]    e_9;
  wire       [1:0]    e_10;
  wire       [1:0]    e_11;
  wire       [1:0]    e_12;
  wire       [1:0]    f_0;
  wire       [1:0]    f_1;
  wire       [1:0]    f_2;
  wire       [1:0]    f_3;
  wire       [1:0]    f_4;
  wire       [1:0]    f_5;
  wire       [1:0]    f_6;
  wire       [1:0]    f_7;
  wire       [1:0]    f_8;
  wire       [1:0]    f_9;
  wire       [1:0]    f_10;
  wire       [1:0]    f_11;
  wire       [1:0]    f_12;
  wire       [1:0]    g_0;
  wire       [1:0]    g_1;
  wire       [1:0]    g_2;
  wire       [1:0]    g_3;
  wire       [1:0]    g_4;
  wire       [1:0]    g_5;
  wire       [1:0]    g_6;
  wire       [1:0]    g_7;
  wire       [1:0]    g_8;
  wire       [1:0]    g_9;
  wire       [1:0]    g_10;
  wire       [1:0]    g_11;
  wire       [1:0]    g_12;
  wire       [1:0]    h_0;
  wire       [1:0]    h_1;
  wire       [1:0]    h_2;
  wire       [1:0]    h_3;
  wire       [1:0]    h_4;
  wire       [1:0]    h_5;
  wire       [1:0]    h_6;
  wire       [1:0]    h_7;
  wire       [1:0]    h_8;
  wire       [1:0]    h_9;
  wire       [1:0]    h_10;
  wire       [1:0]    h_11;
  wire       [1:0]    h_12;
  wire       [1:0]    p_0;
  wire       [1:0]    p_1;
  wire       [1:0]    p_2;
  wire       [1:0]    p_3;
  wire       [1:0]    p_4;
  wire       [1:0]    p_5;
  wire       [1:0]    p_6;
  wire       [1:0]    p_7;
  wire       [1:0]    p_8;
  wire       [1:0]    p_9;
  wire       [1:0]    p_10;
  wire       [1:0]    p_11;
  wire       [1:0]    p_12;
  wire       [1:0]    q_0;
  wire       [1:0]    q_1;
  wire       [1:0]    q_2;
  wire       [1:0]    q_3;
  wire       [1:0]    q_4;
  wire       [1:0]    q_5;
  wire       [1:0]    q_6;
  wire       [1:0]    q_7;
  wire       [1:0]    q_8;
  wire       [1:0]    q_9;
  wire       [1:0]    q_10;
  wire       [1:0]    q_11;
  wire       [1:0]    q_12;

  G4MulTIMaskedN mul1 (
    .io_x_0     (mul1_io_x_0[1:0]   ), //i
    .io_x_1     (mul1_io_x_1[1:0]   ), //i
    .io_x_2     (mul1_io_x_2[1:0]   ), //i
    .io_x_3     (mul1_io_x_3[1:0]   ), //i
    .io_x_4     (mul1_io_x_4[1:0]   ), //i
    .io_x_5     (mul1_io_x_5[1:0]   ), //i
    .io_x_6     (mul1_io_x_6[1:0]   ), //i
    .io_x_7     (mul1_io_x_7[1:0]   ), //i
    .io_x_8     (mul1_io_x_8[1:0]   ), //i
    .io_x_9     (mul1_io_x_9[1:0]   ), //i
    .io_x_10    (mul1_io_x_10[1:0]  ), //i
    .io_x_11    (mul1_io_x_11[1:0]  ), //i
    .io_x_12    (mul1_io_x_12[1:0]  ), //i
    .io_y_0     (mul1_io_y_0[1:0]   ), //i
    .io_y_1     (mul1_io_y_1[1:0]   ), //i
    .io_y_2     (mul1_io_y_2[1:0]   ), //i
    .io_y_3     (mul1_io_y_3[1:0]   ), //i
    .io_y_4     (mul1_io_y_4[1:0]   ), //i
    .io_y_5     (mul1_io_y_5[1:0]   ), //i
    .io_y_6     (mul1_io_y_6[1:0]   ), //i
    .io_y_7     (mul1_io_y_7[1:0]   ), //i
    .io_y_8     (mul1_io_y_8[1:0]   ), //i
    .io_y_9     (mul1_io_y_9[1:0]   ), //i
    .io_y_10    (mul1_io_y_10[1:0]  ), //i
    .io_y_11    (mul1_io_y_11[1:0]  ), //i
    .io_y_12    (mul1_io_y_12[1:0]  ), //i
    .io_z_0     (mul1_io_z_0[1:0]   ), //o
    .io_z_1     (mul1_io_z_1[1:0]   ), //o
    .io_z_2     (mul1_io_z_2[1:0]   ), //o
    .io_z_3     (mul1_io_z_3[1:0]   ), //o
    .io_z_4     (mul1_io_z_4[1:0]   ), //o
    .io_z_5     (mul1_io_z_5[1:0]   ), //o
    .io_z_6     (mul1_io_z_6[1:0]   ), //o
    .io_z_7     (mul1_io_z_7[1:0]   ), //o
    .io_z_8     (mul1_io_z_8[1:0]   ), //o
    .io_z_9     (mul1_io_z_9[1:0]   ), //o
    .io_z_10    (mul1_io_z_10[1:0]  ), //o
    .io_z_11    (mul1_io_z_11[1:0]  ), //o
    .io_z_12    (mul1_io_z_12[1:0]  ), //o
    .clk        (clk                ), //i
    .reset      (reset              )  //i
  );
  G4MulTIMaskedN mul2 (
    .io_x_0     (a_0[1:0]           ), //i
    .io_x_1     (a_1[1:0]           ), //i
    .io_x_2     (a_2[1:0]           ), //i
    .io_x_3     (a_3[1:0]           ), //i
    .io_x_4     (a_4[1:0]           ), //i
    .io_x_5     (a_5[1:0]           ), //i
    .io_x_6     (a_6[1:0]           ), //i
    .io_x_7     (a_7[1:0]           ), //i
    .io_x_8     (a_8[1:0]           ), //i
    .io_x_9     (a_9[1:0]           ), //i
    .io_x_10    (a_10[1:0]          ), //i
    .io_x_11    (a_11[1:0]          ), //i
    .io_x_12    (a_12[1:0]          ), //i
    .io_y_0     (c_0[1:0]           ), //i
    .io_y_1     (c_1[1:0]           ), //i
    .io_y_2     (c_2[1:0]           ), //i
    .io_y_3     (c_3[1:0]           ), //i
    .io_y_4     (c_4[1:0]           ), //i
    .io_y_5     (c_5[1:0]           ), //i
    .io_y_6     (c_6[1:0]           ), //i
    .io_y_7     (c_7[1:0]           ), //i
    .io_y_8     (c_8[1:0]           ), //i
    .io_y_9     (c_9[1:0]           ), //i
    .io_y_10    (c_10[1:0]          ), //i
    .io_y_11    (c_11[1:0]          ), //i
    .io_y_12    (c_12[1:0]          ), //i
    .io_z_0     (mul2_io_z_0[1:0]   ), //o
    .io_z_1     (mul2_io_z_1[1:0]   ), //o
    .io_z_2     (mul2_io_z_2[1:0]   ), //o
    .io_z_3     (mul2_io_z_3[1:0]   ), //o
    .io_z_4     (mul2_io_z_4[1:0]   ), //o
    .io_z_5     (mul2_io_z_5[1:0]   ), //o
    .io_z_6     (mul2_io_z_6[1:0]   ), //o
    .io_z_7     (mul2_io_z_7[1:0]   ), //o
    .io_z_8     (mul2_io_z_8[1:0]   ), //o
    .io_z_9     (mul2_io_z_9[1:0]   ), //o
    .io_z_10    (mul2_io_z_10[1:0]  ), //o
    .io_z_11    (mul2_io_z_11[1:0]  ), //o
    .io_z_12    (mul2_io_z_12[1:0]  ), //o
    .clk        (clk                ), //i
    .reset      (reset              )  //i
  );
  G4MulTIMaskedN mul3 (
    .io_x_0     (b_0[1:0]           ), //i
    .io_x_1     (b_1[1:0]           ), //i
    .io_x_2     (b_2[1:0]           ), //i
    .io_x_3     (b_3[1:0]           ), //i
    .io_x_4     (b_4[1:0]           ), //i
    .io_x_5     (b_5[1:0]           ), //i
    .io_x_6     (b_6[1:0]           ), //i
    .io_x_7     (b_7[1:0]           ), //i
    .io_x_8     (b_8[1:0]           ), //i
    .io_x_9     (b_9[1:0]           ), //i
    .io_x_10    (b_10[1:0]          ), //i
    .io_x_11    (b_11[1:0]          ), //i
    .io_x_12    (b_12[1:0]          ), //i
    .io_y_0     (d_0[1:0]           ), //i
    .io_y_1     (d_1[1:0]           ), //i
    .io_y_2     (d_2[1:0]           ), //i
    .io_y_3     (d_3[1:0]           ), //i
    .io_y_4     (d_4[1:0]           ), //i
    .io_y_5     (d_5[1:0]           ), //i
    .io_y_6     (d_6[1:0]           ), //i
    .io_y_7     (d_7[1:0]           ), //i
    .io_y_8     (d_8[1:0]           ), //i
    .io_y_9     (d_9[1:0]           ), //i
    .io_y_10    (d_10[1:0]          ), //i
    .io_y_11    (d_11[1:0]          ), //i
    .io_y_12    (d_12[1:0]          ), //i
    .io_z_0     (mul3_io_z_0[1:0]   ), //o
    .io_z_1     (mul3_io_z_1[1:0]   ), //o
    .io_z_2     (mul3_io_z_2[1:0]   ), //o
    .io_z_3     (mul3_io_z_3[1:0]   ), //o
    .io_z_4     (mul3_io_z_4[1:0]   ), //o
    .io_z_5     (mul3_io_z_5[1:0]   ), //o
    .io_z_6     (mul3_io_z_6[1:0]   ), //o
    .io_z_7     (mul3_io_z_7[1:0]   ), //o
    .io_z_8     (mul3_io_z_8[1:0]   ), //o
    .io_z_9     (mul3_io_z_9[1:0]   ), //o
    .io_z_10    (mul3_io_z_10[1:0]  ), //o
    .io_z_11    (mul3_io_z_11[1:0]  ), //o
    .io_z_12    (mul3_io_z_12[1:0]  ), //o
    .clk        (clk                ), //i
    .reset      (reset              )  //i
  );
  G4ScaleN g4ScaleN_52 (
    .io_t    (e_0[1:0]               ), //i
    .io_x    (g4ScaleN_52_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_53 (
    .io_t    (e_1[1:0]               ), //i
    .io_x    (g4ScaleN_53_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_54 (
    .io_t    (e_2[1:0]               ), //i
    .io_x    (g4ScaleN_54_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_55 (
    .io_t    (e_3[1:0]               ), //i
    .io_x    (g4ScaleN_55_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_56 (
    .io_t    (e_4[1:0]               ), //i
    .io_x    (g4ScaleN_56_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_57 (
    .io_t    (e_5[1:0]               ), //i
    .io_x    (g4ScaleN_57_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_58 (
    .io_t    (e_6[1:0]               ), //i
    .io_x    (g4ScaleN_58_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_59 (
    .io_t    (e_7[1:0]               ), //i
    .io_x    (g4ScaleN_59_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_60 (
    .io_t    (e_8[1:0]               ), //i
    .io_x    (g4ScaleN_60_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_61 (
    .io_t    (e_9[1:0]               ), //i
    .io_x    (g4ScaleN_61_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_62 (
    .io_t    (e_10[1:0]              ), //i
    .io_x    (g4ScaleN_62_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_63 (
    .io_t    (e_11[1:0]              ), //i
    .io_x    (g4ScaleN_63_io_x[1:0]  )  //o
  );
  G4ScaleN g4ScaleN_64 (
    .io_t    (e_12[1:0]              ), //i
    .io_x    (g4ScaleN_64_io_x[1:0]  )  //o
  );
  assign dummy = 1'b0;
  assign a_0 = io_x_0[3 : 2];
  assign b_0 = io_x_0[1 : 0];
  assign c_0 = io_y_0[3 : 2];
  assign d_0 = io_y_0[1 : 0];
  assign a_1 = io_x_1[3 : 2];
  assign b_1 = io_x_1[1 : 0];
  assign c_1 = io_y_1[3 : 2];
  assign d_1 = io_y_1[1 : 0];
  assign a_2 = io_x_2[3 : 2];
  assign b_2 = io_x_2[1 : 0];
  assign c_2 = io_y_2[3 : 2];
  assign d_2 = io_y_2[1 : 0];
  assign a_3 = io_x_3[3 : 2];
  assign b_3 = io_x_3[1 : 0];
  assign c_3 = io_y_3[3 : 2];
  assign d_3 = io_y_3[1 : 0];
  assign a_4 = io_x_4[3 : 2];
  assign b_4 = io_x_4[1 : 0];
  assign c_4 = io_y_4[3 : 2];
  assign d_4 = io_y_4[1 : 0];
  assign a_5 = io_x_5[3 : 2];
  assign b_5 = io_x_5[1 : 0];
  assign c_5 = io_y_5[3 : 2];
  assign d_5 = io_y_5[1 : 0];
  assign a_6 = io_x_6[3 : 2];
  assign b_6 = io_x_6[1 : 0];
  assign c_6 = io_y_6[3 : 2];
  assign d_6 = io_y_6[1 : 0];
  assign a_7 = io_x_7[3 : 2];
  assign b_7 = io_x_7[1 : 0];
  assign c_7 = io_y_7[3 : 2];
  assign d_7 = io_y_7[1 : 0];
  assign a_8 = io_x_8[3 : 2];
  assign b_8 = io_x_8[1 : 0];
  assign c_8 = io_y_8[3 : 2];
  assign d_8 = io_y_8[1 : 0];
  assign a_9 = io_x_9[3 : 2];
  assign b_9 = io_x_9[1 : 0];
  assign c_9 = io_y_9[3 : 2];
  assign d_9 = io_y_9[1 : 0];
  assign a_10 = io_x_10[3 : 2];
  assign b_10 = io_x_10[1 : 0];
  assign c_10 = io_y_10[3 : 2];
  assign d_10 = io_y_10[1 : 0];
  assign a_11 = io_x_11[3 : 2];
  assign b_11 = io_x_11[1 : 0];
  assign c_11 = io_y_11[3 : 2];
  assign d_11 = io_y_11[1 : 0];
  assign a_12 = io_x_12[3 : 2];
  assign b_12 = io_x_12[1 : 0];
  assign c_12 = io_y_12[3 : 2];
  assign d_12 = io_y_12[1 : 0];
  assign mul1_io_x_0 = (a_0 ^ b_0);
  assign mul1_io_x_1 = (a_1 ^ b_1);
  assign mul1_io_x_2 = (a_2 ^ b_2);
  assign mul1_io_x_3 = (a_3 ^ b_3);
  assign mul1_io_x_4 = (a_4 ^ b_4);
  assign mul1_io_x_5 = (a_5 ^ b_5);
  assign mul1_io_x_6 = (a_6 ^ b_6);
  assign mul1_io_x_7 = (a_7 ^ b_7);
  assign mul1_io_x_8 = (a_8 ^ b_8);
  assign mul1_io_x_9 = (a_9 ^ b_9);
  assign mul1_io_x_10 = (a_10 ^ b_10);
  assign mul1_io_x_11 = (a_11 ^ b_11);
  assign mul1_io_x_12 = (a_12 ^ b_12);
  assign mul1_io_y_0 = (c_0 ^ d_0);
  assign mul1_io_y_1 = (c_1 ^ d_1);
  assign mul1_io_y_2 = (c_2 ^ d_2);
  assign mul1_io_y_3 = (c_3 ^ d_3);
  assign mul1_io_y_4 = (c_4 ^ d_4);
  assign mul1_io_y_5 = (c_5 ^ d_5);
  assign mul1_io_y_6 = (c_6 ^ d_6);
  assign mul1_io_y_7 = (c_7 ^ d_7);
  assign mul1_io_y_8 = (c_8 ^ d_8);
  assign mul1_io_y_9 = (c_9 ^ d_9);
  assign mul1_io_y_10 = (c_10 ^ d_10);
  assign mul1_io_y_11 = (c_11 ^ d_11);
  assign mul1_io_y_12 = (c_12 ^ d_12);
  assign e_0 = mul1_io_z_0;
  assign e_1 = mul1_io_z_1;
  assign e_2 = mul1_io_z_2;
  assign e_3 = mul1_io_z_3;
  assign e_4 = mul1_io_z_4;
  assign e_5 = mul1_io_z_5;
  assign e_6 = mul1_io_z_6;
  assign e_7 = mul1_io_z_7;
  assign e_8 = mul1_io_z_8;
  assign e_9 = mul1_io_z_9;
  assign e_10 = mul1_io_z_10;
  assign e_11 = mul1_io_z_11;
  assign e_12 = mul1_io_z_12;
  assign f_0 = g4ScaleN_52_io_x;
  assign f_1 = g4ScaleN_53_io_x;
  assign f_2 = g4ScaleN_54_io_x;
  assign f_3 = g4ScaleN_55_io_x;
  assign f_4 = g4ScaleN_56_io_x;
  assign f_5 = g4ScaleN_57_io_x;
  assign f_6 = g4ScaleN_58_io_x;
  assign f_7 = g4ScaleN_59_io_x;
  assign f_8 = g4ScaleN_60_io_x;
  assign f_9 = g4ScaleN_61_io_x;
  assign f_10 = g4ScaleN_62_io_x;
  assign f_11 = g4ScaleN_63_io_x;
  assign f_12 = g4ScaleN_64_io_x;
  assign g_0 = mul2_io_z_0;
  assign g_1 = mul2_io_z_1;
  assign g_2 = mul2_io_z_2;
  assign g_3 = mul2_io_z_3;
  assign g_4 = mul2_io_z_4;
  assign g_5 = mul2_io_z_5;
  assign g_6 = mul2_io_z_6;
  assign g_7 = mul2_io_z_7;
  assign g_8 = mul2_io_z_8;
  assign g_9 = mul2_io_z_9;
  assign g_10 = mul2_io_z_10;
  assign g_11 = mul2_io_z_11;
  assign g_12 = mul2_io_z_12;
  assign h_0 = mul3_io_z_0;
  assign h_1 = mul3_io_z_1;
  assign h_2 = mul3_io_z_2;
  assign h_3 = mul3_io_z_3;
  assign h_4 = mul3_io_z_4;
  assign h_5 = mul3_io_z_5;
  assign h_6 = mul3_io_z_6;
  assign h_7 = mul3_io_z_7;
  assign h_8 = mul3_io_z_8;
  assign h_9 = mul3_io_z_9;
  assign h_10 = mul3_io_z_10;
  assign h_11 = mul3_io_z_11;
  assign h_12 = mul3_io_z_12;
  assign p_0 = (f_0 ^ g_0);
  assign p_1 = (f_1 ^ g_1);
  assign p_2 = (f_2 ^ g_2);
  assign p_3 = (f_3 ^ g_3);
  assign p_4 = (f_4 ^ g_4);
  assign p_5 = (f_5 ^ g_5);
  assign p_6 = (f_6 ^ g_6);
  assign p_7 = (f_7 ^ g_7);
  assign p_8 = (f_8 ^ g_8);
  assign p_9 = (f_9 ^ g_9);
  assign p_10 = (f_10 ^ g_10);
  assign p_11 = (f_11 ^ g_11);
  assign p_12 = (f_12 ^ g_12);
  assign q_0 = (f_0 ^ h_0);
  assign q_1 = (f_1 ^ h_1);
  assign q_2 = (f_2 ^ h_2);
  assign q_3 = (f_3 ^ h_3);
  assign q_4 = (f_4 ^ h_4);
  assign q_5 = (f_5 ^ h_5);
  assign q_6 = (f_6 ^ h_6);
  assign q_7 = (f_7 ^ h_7);
  assign q_8 = (f_8 ^ h_8);
  assign q_9 = (f_9 ^ h_9);
  assign q_10 = (f_10 ^ h_10);
  assign q_11 = (f_11 ^ h_11);
  assign q_12 = (f_12 ^ h_12);
  assign io_z_0 = {p_0,q_0};
  assign io_z_1 = {p_1,q_1};
  assign io_z_2 = {p_2,q_2};
  assign io_z_3 = {p_3,q_3};
  assign io_z_4 = {p_4,q_4};
  assign io_z_5 = {p_5,q_5};
  assign io_z_6 = {p_6,q_6};
  assign io_z_7 = {p_7,q_7};
  assign io_z_8 = {p_8,q_8};
  assign io_z_9 = {p_9,q_9};
  assign io_z_10 = {p_10,q_10};
  assign io_z_11 = {p_11,q_11};
  assign io_z_12 = {p_12,q_12};

endmodule

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN2 replaced by G4ScaleN2

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

module G4ScaleN2 (
  input      [1:0]    io_t,
  output     [1:0]    io_x
);


  assign io_x = {(io_t[1] ^ io_t[0]),io_t[1]};

endmodule

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

//G4Sq replaced by G4Sq

//G4ScaleN replaced by G4ScaleN

module G4Sq (
  input      [1:0]    io_t,
  output     [1:0]    io_x
);


  assign io_x = {io_t[0],io_t[1]};

endmodule

//G4MulTIMaskedN replaced by G4MulTIMaskedN

//G4MulTIMaskedN replaced by G4MulTIMaskedN

//G4MulTIMaskedN replaced by G4MulTIMaskedN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4MulTIMaskedN replaced by G4MulTIMaskedN

//G4MulTIMaskedN replaced by G4MulTIMaskedN

//G4MulTIMaskedN replaced by G4MulTIMaskedN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4MulTIMaskedN replaced by G4MulTIMaskedN

//G4MulTIMaskedN replaced by G4MulTIMaskedN

//G4MulTIMaskedN replaced by G4MulTIMaskedN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

//G4ScaleN replaced by G4ScaleN

module G4ScaleN (
  input      [1:0]    io_t,
  output     [1:0]    io_x
);


  assign io_x = {io_t[0],(io_t[1] ^ io_t[0])};

endmodule

//G4MulTIMaskedN replaced by G4MulTIMaskedN

//G4MulTIMaskedN replaced by G4MulTIMaskedN

module G4MulTIMaskedN (
  input      [1:0]    io_x_0,
  input      [1:0]    io_x_1,
  input      [1:0]    io_x_2,
  input      [1:0]    io_x_3,
  input      [1:0]    io_x_4,
  input      [1:0]    io_x_5,
  input      [1:0]    io_x_6,
  input      [1:0]    io_x_7,
  input      [1:0]    io_x_8,
  input      [1:0]    io_x_9,
  input      [1:0]    io_x_10,
  input      [1:0]    io_x_11,
  input      [1:0]    io_x_12,
  input      [1:0]    io_y_0,
  input      [1:0]    io_y_1,
  input      [1:0]    io_y_2,
  input      [1:0]    io_y_3,
  input      [1:0]    io_y_4,
  input      [1:0]    io_y_5,
  input      [1:0]    io_y_6,
  input      [1:0]    io_y_7,
  input      [1:0]    io_y_8,
  input      [1:0]    io_y_9,
  input      [1:0]    io_y_10,
  input      [1:0]    io_y_11,
  input      [1:0]    io_y_12,
  output     [1:0]    io_z_0,
  output     [1:0]    io_z_1,
  output     [1:0]    io_z_2,
  output     [1:0]    io_z_3,
  output     [1:0]    io_z_4,
  output     [1:0]    io_z_5,
  output     [1:0]    io_z_6,
  output     [1:0]    io_z_7,
  output     [1:0]    io_z_8,
  output     [1:0]    io_z_9,
  output     [1:0]    io_z_10,
  output     [1:0]    io_z_11,
  output     [1:0]    io_z_12,
  input               clk,
  input               reset
);

  wire                dummy;
  wire                a_0;
  wire                a_1;
  wire                a_2;
  wire                a_3;
  wire                a_4;
  wire                a_5;
  wire                a_6;
  wire                a_7;
  wire                a_8;
  wire                a_9;
  wire                a_10;
  wire                a_11;
  wire                a_12;
  wire                b_0;
  wire                b_1;
  wire                b_2;
  wire                b_3;
  wire                b_4;
  wire                b_5;
  wire                b_6;
  wire                b_7;
  wire                b_8;
  wire                b_9;
  wire                b_10;
  wire                b_11;
  wire                b_12;
  wire                c_0;
  wire                c_1;
  wire                c_2;
  wire                c_3;
  wire                c_4;
  wire                c_5;
  wire                c_6;
  wire                c_7;
  wire                c_8;
  wire                c_9;
  wire                c_10;
  wire                c_11;
  wire                c_12;
  wire                d_0;
  wire                d_1;
  wire                d_2;
  wire                d_3;
  wire                d_4;
  wire                d_5;
  wire                d_6;
  wire                d_7;
  wire                d_8;
  wire                d_9;
  wire                d_10;
  wire                d_11;
  wire                d_12;
  reg        [12:0]   e_0;
  reg        [12:0]   e_1;
  reg        [12:0]   e_2;
  reg        [12:0]   e_3;
  reg        [12:0]   e_4;
  reg        [12:0]   e_5;
  reg        [12:0]   e_6;
  reg        [12:0]   e_7;
  reg        [12:0]   e_8;
  reg        [12:0]   e_9;
  reg        [12:0]   e_10;
  reg        [12:0]   e_11;
  reg        [12:0]   e_12;
  reg        [12:0]   f_0;
  reg        [12:0]   f_1;
  reg        [12:0]   f_2;
  reg        [12:0]   f_3;
  reg        [12:0]   f_4;
  reg        [12:0]   f_5;
  reg        [12:0]   f_6;
  reg        [12:0]   f_7;
  reg        [12:0]   f_8;
  reg        [12:0]   f_9;
  reg        [12:0]   f_10;
  reg        [12:0]   f_11;
  reg        [12:0]   f_12;
  wire                ac_0;
  wire                ac_1;
  wire                ac_2;
  wire                ac_3;
  wire                ac_4;
  wire                ac_5;
  wire                ac_6;
  wire                ac_7;
  wire                ac_8;
  wire                ac_9;
  wire                ac_10;
  wire                ac_11;
  wire                ac_12;
  wire                ac_13;
  wire                ac_14;
  wire                ac_15;
  wire                ac_16;
  wire                ac_17;
  wire                ac_18;
  wire                ac_19;
  wire                ac_20;
  wire                ac_21;
  wire                ac_22;
  wire                ac_23;
  wire                ac_24;
  wire                ac_25;
  wire                ac_26;
  wire                ac_27;
  wire                ac_28;
  wire                ac_29;
  wire                ac_30;
  wire                ac_31;
  wire                ac_32;
  wire                ac_33;
  wire                ac_34;
  wire                ac_35;
  wire                ac_36;
  wire                ac_37;
  wire                ac_38;
  wire                ac_39;
  wire                ac_40;
  wire                ac_41;
  wire                ac_42;
  wire                ac_43;
  wire                ac_44;
  wire                ac_45;
  wire                ac_46;
  wire                ac_47;
  wire                ac_48;
  wire                ac_49;
  wire                ac_50;
  wire                ac_51;
  wire                ac_52;
  wire                ac_53;
  wire                ac_54;
  wire                ac_55;
  wire                ac_56;
  wire                ac_57;
  wire                ac_58;
  wire                ac_59;
  wire                ac_60;
  wire                ac_61;
  wire                ac_62;
  wire                ac_63;
  wire                ac_64;
  wire                ac_65;
  wire                ac_66;
  wire                ac_67;
  wire                ac_68;
  wire                ac_69;
  wire                ac_70;
  wire                ac_71;
  wire                ac_72;
  wire                ac_73;
  wire                ac_74;
  wire                ac_75;
  wire                ac_76;
  wire                ac_77;
  wire                ac_78;
  wire                ac_79;
  wire                ac_80;
  wire                ac_81;
  wire                ac_82;
  wire                ac_83;
  wire                ac_84;
  wire                ac_85;
  wire                ac_86;
  wire                ac_87;
  wire                ac_88;
  wire                ac_89;
  wire                ac_90;
  wire                ac_91;
  wire                ac_92;
  wire                ac_93;
  wire                ac_94;
  wire                ac_95;
  wire                ac_96;
  wire                ac_97;
  wire                ac_98;
  wire                ac_99;
  wire                ac_100;
  wire                ac_101;
  wire                ac_102;
  wire                ac_103;
  wire                ac_104;
  wire                ac_105;
  wire                ac_106;
  wire                ac_107;
  wire                ac_108;
  wire                ac_109;
  wire                ac_110;
  wire                ac_111;
  wire                ac_112;
  wire                ac_113;
  wire                ac_114;
  wire                ac_115;
  wire                ac_116;
  wire                ac_117;
  wire                ac_118;
  wire                ac_119;
  wire                ac_120;
  wire                ac_121;
  wire                ac_122;
  wire                ac_123;
  wire                ac_124;
  wire                ac_125;
  wire                ac_126;
  wire                ac_127;
  wire                ac_128;
  wire                ac_129;
  wire                ac_130;
  wire                ac_131;
  wire                ac_132;
  wire                ac_133;
  wire                ac_134;
  wire                ac_135;
  wire                ac_136;
  wire                ac_137;
  wire                ac_138;
  wire                ac_139;
  wire                ac_140;
  wire                ac_141;
  wire                ac_142;
  wire                ac_143;
  wire                ac_144;
  wire                ac_145;
  wire                ac_146;
  wire                ac_147;
  wire                ac_148;
  wire                ac_149;
  wire                ac_150;
  wire                ac_151;
  wire                ac_152;
  wire                ac_153;
  wire                ac_154;
  wire                ac_155;
  wire                ac_156;
  wire                ac_157;
  wire                ac_158;
  wire                ac_159;
  wire                ac_160;
  wire                ac_161;
  wire                ac_162;
  wire                ac_163;
  wire                ac_164;
  wire                ac_165;
  wire                ac_166;
  wire                ac_167;
  wire                ac_168;
  wire                ad_0;
  wire                ad_1;
  wire                ad_2;
  wire                ad_3;
  wire                ad_4;
  wire                ad_5;
  wire                ad_6;
  wire                ad_7;
  wire                ad_8;
  wire                ad_9;
  wire                ad_10;
  wire                ad_11;
  wire                ad_12;
  wire                ad_13;
  wire                ad_14;
  wire                ad_15;
  wire                ad_16;
  wire                ad_17;
  wire                ad_18;
  wire                ad_19;
  wire                ad_20;
  wire                ad_21;
  wire                ad_22;
  wire                ad_23;
  wire                ad_24;
  wire                ad_25;
  wire                ad_26;
  wire                ad_27;
  wire                ad_28;
  wire                ad_29;
  wire                ad_30;
  wire                ad_31;
  wire                ad_32;
  wire                ad_33;
  wire                ad_34;
  wire                ad_35;
  wire                ad_36;
  wire                ad_37;
  wire                ad_38;
  wire                ad_39;
  wire                ad_40;
  wire                ad_41;
  wire                ad_42;
  wire                ad_43;
  wire                ad_44;
  wire                ad_45;
  wire                ad_46;
  wire                ad_47;
  wire                ad_48;
  wire                ad_49;
  wire                ad_50;
  wire                ad_51;
  wire                ad_52;
  wire                ad_53;
  wire                ad_54;
  wire                ad_55;
  wire                ad_56;
  wire                ad_57;
  wire                ad_58;
  wire                ad_59;
  wire                ad_60;
  wire                ad_61;
  wire                ad_62;
  wire                ad_63;
  wire                ad_64;
  wire                ad_65;
  wire                ad_66;
  wire                ad_67;
  wire                ad_68;
  wire                ad_69;
  wire                ad_70;
  wire                ad_71;
  wire                ad_72;
  wire                ad_73;
  wire                ad_74;
  wire                ad_75;
  wire                ad_76;
  wire                ad_77;
  wire                ad_78;
  wire                ad_79;
  wire                ad_80;
  wire                ad_81;
  wire                ad_82;
  wire                ad_83;
  wire                ad_84;
  wire                ad_85;
  wire                ad_86;
  wire                ad_87;
  wire                ad_88;
  wire                ad_89;
  wire                ad_90;
  wire                ad_91;
  wire                ad_92;
  wire                ad_93;
  wire                ad_94;
  wire                ad_95;
  wire                ad_96;
  wire                ad_97;
  wire                ad_98;
  wire                ad_99;
  wire                ad_100;
  wire                ad_101;
  wire                ad_102;
  wire                ad_103;
  wire                ad_104;
  wire                ad_105;
  wire                ad_106;
  wire                ad_107;
  wire                ad_108;
  wire                ad_109;
  wire                ad_110;
  wire                ad_111;
  wire                ad_112;
  wire                ad_113;
  wire                ad_114;
  wire                ad_115;
  wire                ad_116;
  wire                ad_117;
  wire                ad_118;
  wire                ad_119;
  wire                ad_120;
  wire                ad_121;
  wire                ad_122;
  wire                ad_123;
  wire                ad_124;
  wire                ad_125;
  wire                ad_126;
  wire                ad_127;
  wire                ad_128;
  wire                ad_129;
  wire                ad_130;
  wire                ad_131;
  wire                ad_132;
  wire                ad_133;
  wire                ad_134;
  wire                ad_135;
  wire                ad_136;
  wire                ad_137;
  wire                ad_138;
  wire                ad_139;
  wire                ad_140;
  wire                ad_141;
  wire                ad_142;
  wire                ad_143;
  wire                ad_144;
  wire                ad_145;
  wire                ad_146;
  wire                ad_147;
  wire                ad_148;
  wire                ad_149;
  wire                ad_150;
  wire                ad_151;
  wire                ad_152;
  wire                ad_153;
  wire                ad_154;
  wire                ad_155;
  wire                ad_156;
  wire                ad_157;
  wire                ad_158;
  wire                ad_159;
  wire                ad_160;
  wire                ad_161;
  wire                ad_162;
  wire                ad_163;
  wire                ad_164;
  wire                ad_165;
  wire                ad_166;
  wire                ad_167;
  wire                ad_168;
  wire                bc_0;
  wire                bc_1;
  wire                bc_2;
  wire                bc_3;
  wire                bc_4;
  wire                bc_5;
  wire                bc_6;
  wire                bc_7;
  wire                bc_8;
  wire                bc_9;
  wire                bc_10;
  wire                bc_11;
  wire                bc_12;
  wire                bc_13;
  wire                bc_14;
  wire                bc_15;
  wire                bc_16;
  wire                bc_17;
  wire                bc_18;
  wire                bc_19;
  wire                bc_20;
  wire                bc_21;
  wire                bc_22;
  wire                bc_23;
  wire                bc_24;
  wire                bc_25;
  wire                bc_26;
  wire                bc_27;
  wire                bc_28;
  wire                bc_29;
  wire                bc_30;
  wire                bc_31;
  wire                bc_32;
  wire                bc_33;
  wire                bc_34;
  wire                bc_35;
  wire                bc_36;
  wire                bc_37;
  wire                bc_38;
  wire                bc_39;
  wire                bc_40;
  wire                bc_41;
  wire                bc_42;
  wire                bc_43;
  wire                bc_44;
  wire                bc_45;
  wire                bc_46;
  wire                bc_47;
  wire                bc_48;
  wire                bc_49;
  wire                bc_50;
  wire                bc_51;
  wire                bc_52;
  wire                bc_53;
  wire                bc_54;
  wire                bc_55;
  wire                bc_56;
  wire                bc_57;
  wire                bc_58;
  wire                bc_59;
  wire                bc_60;
  wire                bc_61;
  wire                bc_62;
  wire                bc_63;
  wire                bc_64;
  wire                bc_65;
  wire                bc_66;
  wire                bc_67;
  wire                bc_68;
  wire                bc_69;
  wire                bc_70;
  wire                bc_71;
  wire                bc_72;
  wire                bc_73;
  wire                bc_74;
  wire                bc_75;
  wire                bc_76;
  wire                bc_77;
  wire                bc_78;
  wire                bc_79;
  wire                bc_80;
  wire                bc_81;
  wire                bc_82;
  wire                bc_83;
  wire                bc_84;
  wire                bc_85;
  wire                bc_86;
  wire                bc_87;
  wire                bc_88;
  wire                bc_89;
  wire                bc_90;
  wire                bc_91;
  wire                bc_92;
  wire                bc_93;
  wire                bc_94;
  wire                bc_95;
  wire                bc_96;
  wire                bc_97;
  wire                bc_98;
  wire                bc_99;
  wire                bc_100;
  wire                bc_101;
  wire                bc_102;
  wire                bc_103;
  wire                bc_104;
  wire                bc_105;
  wire                bc_106;
  wire                bc_107;
  wire                bc_108;
  wire                bc_109;
  wire                bc_110;
  wire                bc_111;
  wire                bc_112;
  wire                bc_113;
  wire                bc_114;
  wire                bc_115;
  wire                bc_116;
  wire                bc_117;
  wire                bc_118;
  wire                bc_119;
  wire                bc_120;
  wire                bc_121;
  wire                bc_122;
  wire                bc_123;
  wire                bc_124;
  wire                bc_125;
  wire                bc_126;
  wire                bc_127;
  wire                bc_128;
  wire                bc_129;
  wire                bc_130;
  wire                bc_131;
  wire                bc_132;
  wire                bc_133;
  wire                bc_134;
  wire                bc_135;
  wire                bc_136;
  wire                bc_137;
  wire                bc_138;
  wire                bc_139;
  wire                bc_140;
  wire                bc_141;
  wire                bc_142;
  wire                bc_143;
  wire                bc_144;
  wire                bc_145;
  wire                bc_146;
  wire                bc_147;
  wire                bc_148;
  wire                bc_149;
  wire                bc_150;
  wire                bc_151;
  wire                bc_152;
  wire                bc_153;
  wire                bc_154;
  wire                bc_155;
  wire                bc_156;
  wire                bc_157;
  wire                bc_158;
  wire                bc_159;
  wire                bc_160;
  wire                bc_161;
  wire                bc_162;
  wire                bc_163;
  wire                bc_164;
  wire                bc_165;
  wire                bc_166;
  wire                bc_167;
  wire                bc_168;
  wire                bd_0;
  wire                bd_1;
  wire                bd_2;
  wire                bd_3;
  wire                bd_4;
  wire                bd_5;
  wire                bd_6;
  wire                bd_7;
  wire                bd_8;
  wire                bd_9;
  wire                bd_10;
  wire                bd_11;
  wire                bd_12;
  wire                bd_13;
  wire                bd_14;
  wire                bd_15;
  wire                bd_16;
  wire                bd_17;
  wire                bd_18;
  wire                bd_19;
  wire                bd_20;
  wire                bd_21;
  wire                bd_22;
  wire                bd_23;
  wire                bd_24;
  wire                bd_25;
  wire                bd_26;
  wire                bd_27;
  wire                bd_28;
  wire                bd_29;
  wire                bd_30;
  wire                bd_31;
  wire                bd_32;
  wire                bd_33;
  wire                bd_34;
  wire                bd_35;
  wire                bd_36;
  wire                bd_37;
  wire                bd_38;
  wire                bd_39;
  wire                bd_40;
  wire                bd_41;
  wire                bd_42;
  wire                bd_43;
  wire                bd_44;
  wire                bd_45;
  wire                bd_46;
  wire                bd_47;
  wire                bd_48;
  wire                bd_49;
  wire                bd_50;
  wire                bd_51;
  wire                bd_52;
  wire                bd_53;
  wire                bd_54;
  wire                bd_55;
  wire                bd_56;
  wire                bd_57;
  wire                bd_58;
  wire                bd_59;
  wire                bd_60;
  wire                bd_61;
  wire                bd_62;
  wire                bd_63;
  wire                bd_64;
  wire                bd_65;
  wire                bd_66;
  wire                bd_67;
  wire                bd_68;
  wire                bd_69;
  wire                bd_70;
  wire                bd_71;
  wire                bd_72;
  wire                bd_73;
  wire                bd_74;
  wire                bd_75;
  wire                bd_76;
  wire                bd_77;
  wire                bd_78;
  wire                bd_79;
  wire                bd_80;
  wire                bd_81;
  wire                bd_82;
  wire                bd_83;
  wire                bd_84;
  wire                bd_85;
  wire                bd_86;
  wire                bd_87;
  wire                bd_88;
  wire                bd_89;
  wire                bd_90;
  wire                bd_91;
  wire                bd_92;
  wire                bd_93;
  wire                bd_94;
  wire                bd_95;
  wire                bd_96;
  wire                bd_97;
  wire                bd_98;
  wire                bd_99;
  wire                bd_100;
  wire                bd_101;
  wire                bd_102;
  wire                bd_103;
  wire                bd_104;
  wire                bd_105;
  wire                bd_106;
  wire                bd_107;
  wire                bd_108;
  wire                bd_109;
  wire                bd_110;
  wire                bd_111;
  wire                bd_112;
  wire                bd_113;
  wire                bd_114;
  wire                bd_115;
  wire                bd_116;
  wire                bd_117;
  wire                bd_118;
  wire                bd_119;
  wire                bd_120;
  wire                bd_121;
  wire                bd_122;
  wire                bd_123;
  wire                bd_124;
  wire                bd_125;
  wire                bd_126;
  wire                bd_127;
  wire                bd_128;
  wire                bd_129;
  wire                bd_130;
  wire                bd_131;
  wire                bd_132;
  wire                bd_133;
  wire                bd_134;
  wire                bd_135;
  wire                bd_136;
  wire                bd_137;
  wire                bd_138;
  wire                bd_139;
  wire                bd_140;
  wire                bd_141;
  wire                bd_142;
  wire                bd_143;
  wire                bd_144;
  wire                bd_145;
  wire                bd_146;
  wire                bd_147;
  wire                bd_148;
  wire                bd_149;
  wire                bd_150;
  wire                bd_151;
  wire                bd_152;
  wire                bd_153;
  wire                bd_154;
  wire                bd_155;
  wire                bd_156;
  wire                bd_157;
  wire                bd_158;
  wire                bd_159;
  wire                bd_160;
  wire                bd_161;
  wire                bd_162;
  wire                bd_163;
  wire                bd_164;
  wire                bd_165;
  wire                bd_166;
  wire                bd_167;
  wire                bd_168;

  assign dummy = 1'b0;
  assign a_0 = io_x_0[1];
  assign b_0 = io_x_0[0];
  assign c_0 = io_y_0[1];
  assign d_0 = io_y_0[0];
  assign a_1 = io_x_1[1];
  assign b_1 = io_x_1[0];
  assign c_1 = io_y_1[1];
  assign d_1 = io_y_1[0];
  assign a_2 = io_x_2[1];
  assign b_2 = io_x_2[0];
  assign c_2 = io_y_2[1];
  assign d_2 = io_y_2[0];
  assign a_3 = io_x_3[1];
  assign b_3 = io_x_3[0];
  assign c_3 = io_y_3[1];
  assign d_3 = io_y_3[0];
  assign a_4 = io_x_4[1];
  assign b_4 = io_x_4[0];
  assign c_4 = io_y_4[1];
  assign d_4 = io_y_4[0];
  assign a_5 = io_x_5[1];
  assign b_5 = io_x_5[0];
  assign c_5 = io_y_5[1];
  assign d_5 = io_y_5[0];
  assign a_6 = io_x_6[1];
  assign b_6 = io_x_6[0];
  assign c_6 = io_y_6[1];
  assign d_6 = io_y_6[0];
  assign a_7 = io_x_7[1];
  assign b_7 = io_x_7[0];
  assign c_7 = io_y_7[1];
  assign d_7 = io_y_7[0];
  assign a_8 = io_x_8[1];
  assign b_8 = io_x_8[0];
  assign c_8 = io_y_8[1];
  assign d_8 = io_y_8[0];
  assign a_9 = io_x_9[1];
  assign b_9 = io_x_9[0];
  assign c_9 = io_y_9[1];
  assign d_9 = io_y_9[0];
  assign a_10 = io_x_10[1];
  assign b_10 = io_x_10[0];
  assign c_10 = io_y_10[1];
  assign d_10 = io_y_10[0];
  assign a_11 = io_x_11[1];
  assign b_11 = io_x_11[0];
  assign c_11 = io_y_11[1];
  assign d_11 = io_y_11[0];
  assign a_12 = io_x_12[1];
  assign b_12 = io_x_12[0];
  assign c_12 = io_y_12[1];
  assign d_12 = io_y_12[0];
  assign ac_0 = (a_0 && c_0);
  assign ad_0 = (a_0 && d_0);
  assign bc_0 = (b_0 && c_0);
  assign bd_0 = (b_0 && d_0);
  assign ac_1 = (a_0 && c_1);
  assign ad_1 = (a_0 && d_1);
  assign bc_1 = (b_0 && c_1);
  assign bd_1 = (b_0 && d_1);
  assign ac_2 = (a_0 && c_2);
  assign ad_2 = (a_0 && d_2);
  assign bc_2 = (b_0 && c_2);
  assign bd_2 = (b_0 && d_2);
  assign ac_3 = (a_0 && c_3);
  assign ad_3 = (a_0 && d_3);
  assign bc_3 = (b_0 && c_3);
  assign bd_3 = (b_0 && d_3);
  assign ac_4 = (a_0 && c_4);
  assign ad_4 = (a_0 && d_4);
  assign bc_4 = (b_0 && c_4);
  assign bd_4 = (b_0 && d_4);
  assign ac_5 = (a_0 && c_5);
  assign ad_5 = (a_0 && d_5);
  assign bc_5 = (b_0 && c_5);
  assign bd_5 = (b_0 && d_5);
  assign ac_6 = (a_0 && c_6);
  assign ad_6 = (a_0 && d_6);
  assign bc_6 = (b_0 && c_6);
  assign bd_6 = (b_0 && d_6);
  assign ac_7 = (a_0 && c_7);
  assign ad_7 = (a_0 && d_7);
  assign bc_7 = (b_0 && c_7);
  assign bd_7 = (b_0 && d_7);
  assign ac_8 = (a_0 && c_8);
  assign ad_8 = (a_0 && d_8);
  assign bc_8 = (b_0 && c_8);
  assign bd_8 = (b_0 && d_8);
  assign ac_9 = (a_0 && c_9);
  assign ad_9 = (a_0 && d_9);
  assign bc_9 = (b_0 && c_9);
  assign bd_9 = (b_0 && d_9);
  assign ac_10 = (a_0 && c_10);
  assign ad_10 = (a_0 && d_10);
  assign bc_10 = (b_0 && c_10);
  assign bd_10 = (b_0 && d_10);
  assign ac_11 = (a_0 && c_11);
  assign ad_11 = (a_0 && d_11);
  assign bc_11 = (b_0 && c_11);
  assign bd_11 = (b_0 && d_11);
  assign ac_12 = (a_0 && c_12);
  assign ad_12 = (a_0 && d_12);
  assign bc_12 = (b_0 && c_12);
  assign bd_12 = (b_0 && d_12);
  assign ac_13 = (a_1 && c_0);
  assign ad_13 = (a_1 && d_0);
  assign bc_13 = (b_1 && c_0);
  assign bd_13 = (b_1 && d_0);
  assign ac_14 = (a_1 && c_1);
  assign ad_14 = (a_1 && d_1);
  assign bc_14 = (b_1 && c_1);
  assign bd_14 = (b_1 && d_1);
  assign ac_15 = (a_1 && c_2);
  assign ad_15 = (a_1 && d_2);
  assign bc_15 = (b_1 && c_2);
  assign bd_15 = (b_1 && d_2);
  assign ac_16 = (a_1 && c_3);
  assign ad_16 = (a_1 && d_3);
  assign bc_16 = (b_1 && c_3);
  assign bd_16 = (b_1 && d_3);
  assign ac_17 = (a_1 && c_4);
  assign ad_17 = (a_1 && d_4);
  assign bc_17 = (b_1 && c_4);
  assign bd_17 = (b_1 && d_4);
  assign ac_18 = (a_1 && c_5);
  assign ad_18 = (a_1 && d_5);
  assign bc_18 = (b_1 && c_5);
  assign bd_18 = (b_1 && d_5);
  assign ac_19 = (a_1 && c_6);
  assign ad_19 = (a_1 && d_6);
  assign bc_19 = (b_1 && c_6);
  assign bd_19 = (b_1 && d_6);
  assign ac_20 = (a_1 && c_7);
  assign ad_20 = (a_1 && d_7);
  assign bc_20 = (b_1 && c_7);
  assign bd_20 = (b_1 && d_7);
  assign ac_21 = (a_1 && c_8);
  assign ad_21 = (a_1 && d_8);
  assign bc_21 = (b_1 && c_8);
  assign bd_21 = (b_1 && d_8);
  assign ac_22 = (a_1 && c_9);
  assign ad_22 = (a_1 && d_9);
  assign bc_22 = (b_1 && c_9);
  assign bd_22 = (b_1 && d_9);
  assign ac_23 = (a_1 && c_10);
  assign ad_23 = (a_1 && d_10);
  assign bc_23 = (b_1 && c_10);
  assign bd_23 = (b_1 && d_10);
  assign ac_24 = (a_1 && c_11);
  assign ad_24 = (a_1 && d_11);
  assign bc_24 = (b_1 && c_11);
  assign bd_24 = (b_1 && d_11);
  assign ac_25 = (a_1 && c_12);
  assign ad_25 = (a_1 && d_12);
  assign bc_25 = (b_1 && c_12);
  assign bd_25 = (b_1 && d_12);
  assign ac_26 = (a_2 && c_0);
  assign ad_26 = (a_2 && d_0);
  assign bc_26 = (b_2 && c_0);
  assign bd_26 = (b_2 && d_0);
  assign ac_27 = (a_2 && c_1);
  assign ad_27 = (a_2 && d_1);
  assign bc_27 = (b_2 && c_1);
  assign bd_27 = (b_2 && d_1);
  assign ac_28 = (a_2 && c_2);
  assign ad_28 = (a_2 && d_2);
  assign bc_28 = (b_2 && c_2);
  assign bd_28 = (b_2 && d_2);
  assign ac_29 = (a_2 && c_3);
  assign ad_29 = (a_2 && d_3);
  assign bc_29 = (b_2 && c_3);
  assign bd_29 = (b_2 && d_3);
  assign ac_30 = (a_2 && c_4);
  assign ad_30 = (a_2 && d_4);
  assign bc_30 = (b_2 && c_4);
  assign bd_30 = (b_2 && d_4);
  assign ac_31 = (a_2 && c_5);
  assign ad_31 = (a_2 && d_5);
  assign bc_31 = (b_2 && c_5);
  assign bd_31 = (b_2 && d_5);
  assign ac_32 = (a_2 && c_6);
  assign ad_32 = (a_2 && d_6);
  assign bc_32 = (b_2 && c_6);
  assign bd_32 = (b_2 && d_6);
  assign ac_33 = (a_2 && c_7);
  assign ad_33 = (a_2 && d_7);
  assign bc_33 = (b_2 && c_7);
  assign bd_33 = (b_2 && d_7);
  assign ac_34 = (a_2 && c_8);
  assign ad_34 = (a_2 && d_8);
  assign bc_34 = (b_2 && c_8);
  assign bd_34 = (b_2 && d_8);
  assign ac_35 = (a_2 && c_9);
  assign ad_35 = (a_2 && d_9);
  assign bc_35 = (b_2 && c_9);
  assign bd_35 = (b_2 && d_9);
  assign ac_36 = (a_2 && c_10);
  assign ad_36 = (a_2 && d_10);
  assign bc_36 = (b_2 && c_10);
  assign bd_36 = (b_2 && d_10);
  assign ac_37 = (a_2 && c_11);
  assign ad_37 = (a_2 && d_11);
  assign bc_37 = (b_2 && c_11);
  assign bd_37 = (b_2 && d_11);
  assign ac_38 = (a_2 && c_12);
  assign ad_38 = (a_2 && d_12);
  assign bc_38 = (b_2 && c_12);
  assign bd_38 = (b_2 && d_12);
  assign ac_39 = (a_3 && c_0);
  assign ad_39 = (a_3 && d_0);
  assign bc_39 = (b_3 && c_0);
  assign bd_39 = (b_3 && d_0);
  assign ac_40 = (a_3 && c_1);
  assign ad_40 = (a_3 && d_1);
  assign bc_40 = (b_3 && c_1);
  assign bd_40 = (b_3 && d_1);
  assign ac_41 = (a_3 && c_2);
  assign ad_41 = (a_3 && d_2);
  assign bc_41 = (b_3 && c_2);
  assign bd_41 = (b_3 && d_2);
  assign ac_42 = (a_3 && c_3);
  assign ad_42 = (a_3 && d_3);
  assign bc_42 = (b_3 && c_3);
  assign bd_42 = (b_3 && d_3);
  assign ac_43 = (a_3 && c_4);
  assign ad_43 = (a_3 && d_4);
  assign bc_43 = (b_3 && c_4);
  assign bd_43 = (b_3 && d_4);
  assign ac_44 = (a_3 && c_5);
  assign ad_44 = (a_3 && d_5);
  assign bc_44 = (b_3 && c_5);
  assign bd_44 = (b_3 && d_5);
  assign ac_45 = (a_3 && c_6);
  assign ad_45 = (a_3 && d_6);
  assign bc_45 = (b_3 && c_6);
  assign bd_45 = (b_3 && d_6);
  assign ac_46 = (a_3 && c_7);
  assign ad_46 = (a_3 && d_7);
  assign bc_46 = (b_3 && c_7);
  assign bd_46 = (b_3 && d_7);
  assign ac_47 = (a_3 && c_8);
  assign ad_47 = (a_3 && d_8);
  assign bc_47 = (b_3 && c_8);
  assign bd_47 = (b_3 && d_8);
  assign ac_48 = (a_3 && c_9);
  assign ad_48 = (a_3 && d_9);
  assign bc_48 = (b_3 && c_9);
  assign bd_48 = (b_3 && d_9);
  assign ac_49 = (a_3 && c_10);
  assign ad_49 = (a_3 && d_10);
  assign bc_49 = (b_3 && c_10);
  assign bd_49 = (b_3 && d_10);
  assign ac_50 = (a_3 && c_11);
  assign ad_50 = (a_3 && d_11);
  assign bc_50 = (b_3 && c_11);
  assign bd_50 = (b_3 && d_11);
  assign ac_51 = (a_3 && c_12);
  assign ad_51 = (a_3 && d_12);
  assign bc_51 = (b_3 && c_12);
  assign bd_51 = (b_3 && d_12);
  assign ac_52 = (a_4 && c_0);
  assign ad_52 = (a_4 && d_0);
  assign bc_52 = (b_4 && c_0);
  assign bd_52 = (b_4 && d_0);
  assign ac_53 = (a_4 && c_1);
  assign ad_53 = (a_4 && d_1);
  assign bc_53 = (b_4 && c_1);
  assign bd_53 = (b_4 && d_1);
  assign ac_54 = (a_4 && c_2);
  assign ad_54 = (a_4 && d_2);
  assign bc_54 = (b_4 && c_2);
  assign bd_54 = (b_4 && d_2);
  assign ac_55 = (a_4 && c_3);
  assign ad_55 = (a_4 && d_3);
  assign bc_55 = (b_4 && c_3);
  assign bd_55 = (b_4 && d_3);
  assign ac_56 = (a_4 && c_4);
  assign ad_56 = (a_4 && d_4);
  assign bc_56 = (b_4 && c_4);
  assign bd_56 = (b_4 && d_4);
  assign ac_57 = (a_4 && c_5);
  assign ad_57 = (a_4 && d_5);
  assign bc_57 = (b_4 && c_5);
  assign bd_57 = (b_4 && d_5);
  assign ac_58 = (a_4 && c_6);
  assign ad_58 = (a_4 && d_6);
  assign bc_58 = (b_4 && c_6);
  assign bd_58 = (b_4 && d_6);
  assign ac_59 = (a_4 && c_7);
  assign ad_59 = (a_4 && d_7);
  assign bc_59 = (b_4 && c_7);
  assign bd_59 = (b_4 && d_7);
  assign ac_60 = (a_4 && c_8);
  assign ad_60 = (a_4 && d_8);
  assign bc_60 = (b_4 && c_8);
  assign bd_60 = (b_4 && d_8);
  assign ac_61 = (a_4 && c_9);
  assign ad_61 = (a_4 && d_9);
  assign bc_61 = (b_4 && c_9);
  assign bd_61 = (b_4 && d_9);
  assign ac_62 = (a_4 && c_10);
  assign ad_62 = (a_4 && d_10);
  assign bc_62 = (b_4 && c_10);
  assign bd_62 = (b_4 && d_10);
  assign ac_63 = (a_4 && c_11);
  assign ad_63 = (a_4 && d_11);
  assign bc_63 = (b_4 && c_11);
  assign bd_63 = (b_4 && d_11);
  assign ac_64 = (a_4 && c_12);
  assign ad_64 = (a_4 && d_12);
  assign bc_64 = (b_4 && c_12);
  assign bd_64 = (b_4 && d_12);
  assign ac_65 = (a_5 && c_0);
  assign ad_65 = (a_5 && d_0);
  assign bc_65 = (b_5 && c_0);
  assign bd_65 = (b_5 && d_0);
  assign ac_66 = (a_5 && c_1);
  assign ad_66 = (a_5 && d_1);
  assign bc_66 = (b_5 && c_1);
  assign bd_66 = (b_5 && d_1);
  assign ac_67 = (a_5 && c_2);
  assign ad_67 = (a_5 && d_2);
  assign bc_67 = (b_5 && c_2);
  assign bd_67 = (b_5 && d_2);
  assign ac_68 = (a_5 && c_3);
  assign ad_68 = (a_5 && d_3);
  assign bc_68 = (b_5 && c_3);
  assign bd_68 = (b_5 && d_3);
  assign ac_69 = (a_5 && c_4);
  assign ad_69 = (a_5 && d_4);
  assign bc_69 = (b_5 && c_4);
  assign bd_69 = (b_5 && d_4);
  assign ac_70 = (a_5 && c_5);
  assign ad_70 = (a_5 && d_5);
  assign bc_70 = (b_5 && c_5);
  assign bd_70 = (b_5 && d_5);
  assign ac_71 = (a_5 && c_6);
  assign ad_71 = (a_5 && d_6);
  assign bc_71 = (b_5 && c_6);
  assign bd_71 = (b_5 && d_6);
  assign ac_72 = (a_5 && c_7);
  assign ad_72 = (a_5 && d_7);
  assign bc_72 = (b_5 && c_7);
  assign bd_72 = (b_5 && d_7);
  assign ac_73 = (a_5 && c_8);
  assign ad_73 = (a_5 && d_8);
  assign bc_73 = (b_5 && c_8);
  assign bd_73 = (b_5 && d_8);
  assign ac_74 = (a_5 && c_9);
  assign ad_74 = (a_5 && d_9);
  assign bc_74 = (b_5 && c_9);
  assign bd_74 = (b_5 && d_9);
  assign ac_75 = (a_5 && c_10);
  assign ad_75 = (a_5 && d_10);
  assign bc_75 = (b_5 && c_10);
  assign bd_75 = (b_5 && d_10);
  assign ac_76 = (a_5 && c_11);
  assign ad_76 = (a_5 && d_11);
  assign bc_76 = (b_5 && c_11);
  assign bd_76 = (b_5 && d_11);
  assign ac_77 = (a_5 && c_12);
  assign ad_77 = (a_5 && d_12);
  assign bc_77 = (b_5 && c_12);
  assign bd_77 = (b_5 && d_12);
  assign ac_78 = (a_6 && c_0);
  assign ad_78 = (a_6 && d_0);
  assign bc_78 = (b_6 && c_0);
  assign bd_78 = (b_6 && d_0);
  assign ac_79 = (a_6 && c_1);
  assign ad_79 = (a_6 && d_1);
  assign bc_79 = (b_6 && c_1);
  assign bd_79 = (b_6 && d_1);
  assign ac_80 = (a_6 && c_2);
  assign ad_80 = (a_6 && d_2);
  assign bc_80 = (b_6 && c_2);
  assign bd_80 = (b_6 && d_2);
  assign ac_81 = (a_6 && c_3);
  assign ad_81 = (a_6 && d_3);
  assign bc_81 = (b_6 && c_3);
  assign bd_81 = (b_6 && d_3);
  assign ac_82 = (a_6 && c_4);
  assign ad_82 = (a_6 && d_4);
  assign bc_82 = (b_6 && c_4);
  assign bd_82 = (b_6 && d_4);
  assign ac_83 = (a_6 && c_5);
  assign ad_83 = (a_6 && d_5);
  assign bc_83 = (b_6 && c_5);
  assign bd_83 = (b_6 && d_5);
  assign ac_84 = (a_6 && c_6);
  assign ad_84 = (a_6 && d_6);
  assign bc_84 = (b_6 && c_6);
  assign bd_84 = (b_6 && d_6);
  assign ac_85 = (a_6 && c_7);
  assign ad_85 = (a_6 && d_7);
  assign bc_85 = (b_6 && c_7);
  assign bd_85 = (b_6 && d_7);
  assign ac_86 = (a_6 && c_8);
  assign ad_86 = (a_6 && d_8);
  assign bc_86 = (b_6 && c_8);
  assign bd_86 = (b_6 && d_8);
  assign ac_87 = (a_6 && c_9);
  assign ad_87 = (a_6 && d_9);
  assign bc_87 = (b_6 && c_9);
  assign bd_87 = (b_6 && d_9);
  assign ac_88 = (a_6 && c_10);
  assign ad_88 = (a_6 && d_10);
  assign bc_88 = (b_6 && c_10);
  assign bd_88 = (b_6 && d_10);
  assign ac_89 = (a_6 && c_11);
  assign ad_89 = (a_6 && d_11);
  assign bc_89 = (b_6 && c_11);
  assign bd_89 = (b_6 && d_11);
  assign ac_90 = (a_6 && c_12);
  assign ad_90 = (a_6 && d_12);
  assign bc_90 = (b_6 && c_12);
  assign bd_90 = (b_6 && d_12);
  assign ac_91 = (a_7 && c_0);
  assign ad_91 = (a_7 && d_0);
  assign bc_91 = (b_7 && c_0);
  assign bd_91 = (b_7 && d_0);
  assign ac_92 = (a_7 && c_1);
  assign ad_92 = (a_7 && d_1);
  assign bc_92 = (b_7 && c_1);
  assign bd_92 = (b_7 && d_1);
  assign ac_93 = (a_7 && c_2);
  assign ad_93 = (a_7 && d_2);
  assign bc_93 = (b_7 && c_2);
  assign bd_93 = (b_7 && d_2);
  assign ac_94 = (a_7 && c_3);
  assign ad_94 = (a_7 && d_3);
  assign bc_94 = (b_7 && c_3);
  assign bd_94 = (b_7 && d_3);
  assign ac_95 = (a_7 && c_4);
  assign ad_95 = (a_7 && d_4);
  assign bc_95 = (b_7 && c_4);
  assign bd_95 = (b_7 && d_4);
  assign ac_96 = (a_7 && c_5);
  assign ad_96 = (a_7 && d_5);
  assign bc_96 = (b_7 && c_5);
  assign bd_96 = (b_7 && d_5);
  assign ac_97 = (a_7 && c_6);
  assign ad_97 = (a_7 && d_6);
  assign bc_97 = (b_7 && c_6);
  assign bd_97 = (b_7 && d_6);
  assign ac_98 = (a_7 && c_7);
  assign ad_98 = (a_7 && d_7);
  assign bc_98 = (b_7 && c_7);
  assign bd_98 = (b_7 && d_7);
  assign ac_99 = (a_7 && c_8);
  assign ad_99 = (a_7 && d_8);
  assign bc_99 = (b_7 && c_8);
  assign bd_99 = (b_7 && d_8);
  assign ac_100 = (a_7 && c_9);
  assign ad_100 = (a_7 && d_9);
  assign bc_100 = (b_7 && c_9);
  assign bd_100 = (b_7 && d_9);
  assign ac_101 = (a_7 && c_10);
  assign ad_101 = (a_7 && d_10);
  assign bc_101 = (b_7 && c_10);
  assign bd_101 = (b_7 && d_10);
  assign ac_102 = (a_7 && c_11);
  assign ad_102 = (a_7 && d_11);
  assign bc_102 = (b_7 && c_11);
  assign bd_102 = (b_7 && d_11);
  assign ac_103 = (a_7 && c_12);
  assign ad_103 = (a_7 && d_12);
  assign bc_103 = (b_7 && c_12);
  assign bd_103 = (b_7 && d_12);
  assign ac_104 = (a_8 && c_0);
  assign ad_104 = (a_8 && d_0);
  assign bc_104 = (b_8 && c_0);
  assign bd_104 = (b_8 && d_0);
  assign ac_105 = (a_8 && c_1);
  assign ad_105 = (a_8 && d_1);
  assign bc_105 = (b_8 && c_1);
  assign bd_105 = (b_8 && d_1);
  assign ac_106 = (a_8 && c_2);
  assign ad_106 = (a_8 && d_2);
  assign bc_106 = (b_8 && c_2);
  assign bd_106 = (b_8 && d_2);
  assign ac_107 = (a_8 && c_3);
  assign ad_107 = (a_8 && d_3);
  assign bc_107 = (b_8 && c_3);
  assign bd_107 = (b_8 && d_3);
  assign ac_108 = (a_8 && c_4);
  assign ad_108 = (a_8 && d_4);
  assign bc_108 = (b_8 && c_4);
  assign bd_108 = (b_8 && d_4);
  assign ac_109 = (a_8 && c_5);
  assign ad_109 = (a_8 && d_5);
  assign bc_109 = (b_8 && c_5);
  assign bd_109 = (b_8 && d_5);
  assign ac_110 = (a_8 && c_6);
  assign ad_110 = (a_8 && d_6);
  assign bc_110 = (b_8 && c_6);
  assign bd_110 = (b_8 && d_6);
  assign ac_111 = (a_8 && c_7);
  assign ad_111 = (a_8 && d_7);
  assign bc_111 = (b_8 && c_7);
  assign bd_111 = (b_8 && d_7);
  assign ac_112 = (a_8 && c_8);
  assign ad_112 = (a_8 && d_8);
  assign bc_112 = (b_8 && c_8);
  assign bd_112 = (b_8 && d_8);
  assign ac_113 = (a_8 && c_9);
  assign ad_113 = (a_8 && d_9);
  assign bc_113 = (b_8 && c_9);
  assign bd_113 = (b_8 && d_9);
  assign ac_114 = (a_8 && c_10);
  assign ad_114 = (a_8 && d_10);
  assign bc_114 = (b_8 && c_10);
  assign bd_114 = (b_8 && d_10);
  assign ac_115 = (a_8 && c_11);
  assign ad_115 = (a_8 && d_11);
  assign bc_115 = (b_8 && c_11);
  assign bd_115 = (b_8 && d_11);
  assign ac_116 = (a_8 && c_12);
  assign ad_116 = (a_8 && d_12);
  assign bc_116 = (b_8 && c_12);
  assign bd_116 = (b_8 && d_12);
  assign ac_117 = (a_9 && c_0);
  assign ad_117 = (a_9 && d_0);
  assign bc_117 = (b_9 && c_0);
  assign bd_117 = (b_9 && d_0);
  assign ac_118 = (a_9 && c_1);
  assign ad_118 = (a_9 && d_1);
  assign bc_118 = (b_9 && c_1);
  assign bd_118 = (b_9 && d_1);
  assign ac_119 = (a_9 && c_2);
  assign ad_119 = (a_9 && d_2);
  assign bc_119 = (b_9 && c_2);
  assign bd_119 = (b_9 && d_2);
  assign ac_120 = (a_9 && c_3);
  assign ad_120 = (a_9 && d_3);
  assign bc_120 = (b_9 && c_3);
  assign bd_120 = (b_9 && d_3);
  assign ac_121 = (a_9 && c_4);
  assign ad_121 = (a_9 && d_4);
  assign bc_121 = (b_9 && c_4);
  assign bd_121 = (b_9 && d_4);
  assign ac_122 = (a_9 && c_5);
  assign ad_122 = (a_9 && d_5);
  assign bc_122 = (b_9 && c_5);
  assign bd_122 = (b_9 && d_5);
  assign ac_123 = (a_9 && c_6);
  assign ad_123 = (a_9 && d_6);
  assign bc_123 = (b_9 && c_6);
  assign bd_123 = (b_9 && d_6);
  assign ac_124 = (a_9 && c_7);
  assign ad_124 = (a_9 && d_7);
  assign bc_124 = (b_9 && c_7);
  assign bd_124 = (b_9 && d_7);
  assign ac_125 = (a_9 && c_8);
  assign ad_125 = (a_9 && d_8);
  assign bc_125 = (b_9 && c_8);
  assign bd_125 = (b_9 && d_8);
  assign ac_126 = (a_9 && c_9);
  assign ad_126 = (a_9 && d_9);
  assign bc_126 = (b_9 && c_9);
  assign bd_126 = (b_9 && d_9);
  assign ac_127 = (a_9 && c_10);
  assign ad_127 = (a_9 && d_10);
  assign bc_127 = (b_9 && c_10);
  assign bd_127 = (b_9 && d_10);
  assign ac_128 = (a_9 && c_11);
  assign ad_128 = (a_9 && d_11);
  assign bc_128 = (b_9 && c_11);
  assign bd_128 = (b_9 && d_11);
  assign ac_129 = (a_9 && c_12);
  assign ad_129 = (a_9 && d_12);
  assign bc_129 = (b_9 && c_12);
  assign bd_129 = (b_9 && d_12);
  assign ac_130 = (a_10 && c_0);
  assign ad_130 = (a_10 && d_0);
  assign bc_130 = (b_10 && c_0);
  assign bd_130 = (b_10 && d_0);
  assign ac_131 = (a_10 && c_1);
  assign ad_131 = (a_10 && d_1);
  assign bc_131 = (b_10 && c_1);
  assign bd_131 = (b_10 && d_1);
  assign ac_132 = (a_10 && c_2);
  assign ad_132 = (a_10 && d_2);
  assign bc_132 = (b_10 && c_2);
  assign bd_132 = (b_10 && d_2);
  assign ac_133 = (a_10 && c_3);
  assign ad_133 = (a_10 && d_3);
  assign bc_133 = (b_10 && c_3);
  assign bd_133 = (b_10 && d_3);
  assign ac_134 = (a_10 && c_4);
  assign ad_134 = (a_10 && d_4);
  assign bc_134 = (b_10 && c_4);
  assign bd_134 = (b_10 && d_4);
  assign ac_135 = (a_10 && c_5);
  assign ad_135 = (a_10 && d_5);
  assign bc_135 = (b_10 && c_5);
  assign bd_135 = (b_10 && d_5);
  assign ac_136 = (a_10 && c_6);
  assign ad_136 = (a_10 && d_6);
  assign bc_136 = (b_10 && c_6);
  assign bd_136 = (b_10 && d_6);
  assign ac_137 = (a_10 && c_7);
  assign ad_137 = (a_10 && d_7);
  assign bc_137 = (b_10 && c_7);
  assign bd_137 = (b_10 && d_7);
  assign ac_138 = (a_10 && c_8);
  assign ad_138 = (a_10 && d_8);
  assign bc_138 = (b_10 && c_8);
  assign bd_138 = (b_10 && d_8);
  assign ac_139 = (a_10 && c_9);
  assign ad_139 = (a_10 && d_9);
  assign bc_139 = (b_10 && c_9);
  assign bd_139 = (b_10 && d_9);
  assign ac_140 = (a_10 && c_10);
  assign ad_140 = (a_10 && d_10);
  assign bc_140 = (b_10 && c_10);
  assign bd_140 = (b_10 && d_10);
  assign ac_141 = (a_10 && c_11);
  assign ad_141 = (a_10 && d_11);
  assign bc_141 = (b_10 && c_11);
  assign bd_141 = (b_10 && d_11);
  assign ac_142 = (a_10 && c_12);
  assign ad_142 = (a_10 && d_12);
  assign bc_142 = (b_10 && c_12);
  assign bd_142 = (b_10 && d_12);
  assign ac_143 = (a_11 && c_0);
  assign ad_143 = (a_11 && d_0);
  assign bc_143 = (b_11 && c_0);
  assign bd_143 = (b_11 && d_0);
  assign ac_144 = (a_11 && c_1);
  assign ad_144 = (a_11 && d_1);
  assign bc_144 = (b_11 && c_1);
  assign bd_144 = (b_11 && d_1);
  assign ac_145 = (a_11 && c_2);
  assign ad_145 = (a_11 && d_2);
  assign bc_145 = (b_11 && c_2);
  assign bd_145 = (b_11 && d_2);
  assign ac_146 = (a_11 && c_3);
  assign ad_146 = (a_11 && d_3);
  assign bc_146 = (b_11 && c_3);
  assign bd_146 = (b_11 && d_3);
  assign ac_147 = (a_11 && c_4);
  assign ad_147 = (a_11 && d_4);
  assign bc_147 = (b_11 && c_4);
  assign bd_147 = (b_11 && d_4);
  assign ac_148 = (a_11 && c_5);
  assign ad_148 = (a_11 && d_5);
  assign bc_148 = (b_11 && c_5);
  assign bd_148 = (b_11 && d_5);
  assign ac_149 = (a_11 && c_6);
  assign ad_149 = (a_11 && d_6);
  assign bc_149 = (b_11 && c_6);
  assign bd_149 = (b_11 && d_6);
  assign ac_150 = (a_11 && c_7);
  assign ad_150 = (a_11 && d_7);
  assign bc_150 = (b_11 && c_7);
  assign bd_150 = (b_11 && d_7);
  assign ac_151 = (a_11 && c_8);
  assign ad_151 = (a_11 && d_8);
  assign bc_151 = (b_11 && c_8);
  assign bd_151 = (b_11 && d_8);
  assign ac_152 = (a_11 && c_9);
  assign ad_152 = (a_11 && d_9);
  assign bc_152 = (b_11 && c_9);
  assign bd_152 = (b_11 && d_9);
  assign ac_153 = (a_11 && c_10);
  assign ad_153 = (a_11 && d_10);
  assign bc_153 = (b_11 && c_10);
  assign bd_153 = (b_11 && d_10);
  assign ac_154 = (a_11 && c_11);
  assign ad_154 = (a_11 && d_11);
  assign bc_154 = (b_11 && c_11);
  assign bd_154 = (b_11 && d_11);
  assign ac_155 = (a_11 && c_12);
  assign ad_155 = (a_11 && d_12);
  assign bc_155 = (b_11 && c_12);
  assign bd_155 = (b_11 && d_12);
  assign ac_156 = (a_12 && c_0);
  assign ad_156 = (a_12 && d_0);
  assign bc_156 = (b_12 && c_0);
  assign bd_156 = (b_12 && d_0);
  assign ac_157 = (a_12 && c_1);
  assign ad_157 = (a_12 && d_1);
  assign bc_157 = (b_12 && c_1);
  assign bd_157 = (b_12 && d_1);
  assign ac_158 = (a_12 && c_2);
  assign ad_158 = (a_12 && d_2);
  assign bc_158 = (b_12 && c_2);
  assign bd_158 = (b_12 && d_2);
  assign ac_159 = (a_12 && c_3);
  assign ad_159 = (a_12 && d_3);
  assign bc_159 = (b_12 && c_3);
  assign bd_159 = (b_12 && d_3);
  assign ac_160 = (a_12 && c_4);
  assign ad_160 = (a_12 && d_4);
  assign bc_160 = (b_12 && c_4);
  assign bd_160 = (b_12 && d_4);
  assign ac_161 = (a_12 && c_5);
  assign ad_161 = (a_12 && d_5);
  assign bc_161 = (b_12 && c_5);
  assign bd_161 = (b_12 && d_5);
  assign ac_162 = (a_12 && c_6);
  assign ad_162 = (a_12 && d_6);
  assign bc_162 = (b_12 && c_6);
  assign bd_162 = (b_12 && d_6);
  assign ac_163 = (a_12 && c_7);
  assign ad_163 = (a_12 && d_7);
  assign bc_163 = (b_12 && c_7);
  assign bd_163 = (b_12 && d_7);
  assign ac_164 = (a_12 && c_8);
  assign ad_164 = (a_12 && d_8);
  assign bc_164 = (b_12 && c_8);
  assign bd_164 = (b_12 && d_8);
  assign ac_165 = (a_12 && c_9);
  assign ad_165 = (a_12 && d_9);
  assign bc_165 = (b_12 && c_9);
  assign bd_165 = (b_12 && d_9);
  assign ac_166 = (a_12 && c_10);
  assign ad_166 = (a_12 && d_10);
  assign bc_166 = (b_12 && c_10);
  assign bd_166 = (b_12 && d_10);
  assign ac_167 = (a_12 && c_11);
  assign ad_167 = (a_12 && d_11);
  assign bc_167 = (b_12 && c_11);
  assign bd_167 = (b_12 && d_11);
  assign ac_168 = (a_12 && c_12);
  assign ad_168 = (a_12 && d_12);
  assign bc_168 = (b_12 && c_12);
  assign bd_168 = (b_12 && d_12);
  always @(*) begin
    e_0[12] = ((bc_0 ^ ad_0) ^ bd_0);
    e_0[0] = ((bc_14 ^ ad_14) ^ bd_14);
    e_0[1] = ((bc_28 ^ ad_28) ^ bd_28);
    e_0[2] = ((bc_42 ^ ad_42) ^ bd_42);
    e_0[3] = ((bc_56 ^ ad_56) ^ bd_56);
    e_0[4] = ((bc_70 ^ ad_70) ^ bd_70);
    e_0[5] = ((bc_84 ^ ad_84) ^ bd_84);
    e_0[6] = ((bc_98 ^ ad_98) ^ bd_98);
    e_0[7] = ((bc_112 ^ ad_112) ^ bd_112);
    e_0[8] = ((bc_126 ^ ad_126) ^ bd_126);
    e_0[9] = ((bc_140 ^ ad_140) ^ bd_140);
    e_0[10] = ((bc_154 ^ ad_154) ^ bd_154);
    e_0[11] = ((bc_168 ^ ad_168) ^ bd_168);
  end

  always @(*) begin
    f_0[12] = ((bc_0 ^ ad_0) ^ ac_0);
    f_0[0] = ((bc_14 ^ ad_14) ^ ac_14);
    f_0[1] = ((bc_28 ^ ad_28) ^ ac_28);
    f_0[2] = ((bc_42 ^ ad_42) ^ ac_42);
    f_0[3] = ((bc_56 ^ ad_56) ^ ac_56);
    f_0[4] = ((bc_70 ^ ad_70) ^ ac_70);
    f_0[5] = ((bc_84 ^ ad_84) ^ ac_84);
    f_0[6] = ((bc_98 ^ ad_98) ^ ac_98);
    f_0[7] = ((bc_112 ^ ad_112) ^ ac_112);
    f_0[8] = ((bc_126 ^ ad_126) ^ ac_126);
    f_0[9] = ((bc_140 ^ ad_140) ^ ac_140);
    f_0[10] = ((bc_154 ^ ad_154) ^ ac_154);
    f_0[11] = ((bc_168 ^ ad_168) ^ ac_168);
  end

  always @(*) begin
    e_1[0] = (((e_0[0] ^ bc_15) ^ ad_15) ^ bd_15);
    e_1[1] = (((e_0[1] ^ bc_2) ^ ad_2) ^ bd_2);
    e_1[2] = (((e_0[2] ^ bc_1) ^ ad_1) ^ bd_1);
    e_1[3] = (((e_0[3] ^ bc_4) ^ ad_4) ^ bd_4);
    e_1[4] = (((e_0[4] ^ bc_3) ^ ad_3) ^ bd_3);
    e_1[5] = (((e_0[5] ^ bc_6) ^ ad_6) ^ bd_6);
    e_1[6] = (((e_0[6] ^ bc_5) ^ ad_5) ^ bd_5);
    e_1[7] = (((e_0[7] ^ bc_8) ^ ad_8) ^ bd_8);
    e_1[8] = (((e_0[8] ^ bc_7) ^ ad_7) ^ bd_7);
    e_1[9] = (((e_0[9] ^ bc_10) ^ ad_10) ^ bd_10);
    e_1[10] = (((e_0[10] ^ bc_9) ^ ad_9) ^ bd_9);
    e_1[11] = (((e_0[11] ^ bc_12) ^ ad_12) ^ bd_12);
    e_1[12] = (((e_0[12] ^ bc_11) ^ ad_11) ^ bd_11);
  end

  always @(*) begin
    f_1[0] = (((f_0[0] ^ bc_15) ^ ad_15) ^ ac_15);
    f_1[1] = (((f_0[1] ^ bc_2) ^ ad_2) ^ ac_2);
    f_1[2] = (((f_0[2] ^ bc_1) ^ ad_1) ^ ac_1);
    f_1[3] = (((f_0[3] ^ bc_4) ^ ad_4) ^ ac_4);
    f_1[4] = (((f_0[4] ^ bc_3) ^ ad_3) ^ ac_3);
    f_1[5] = (((f_0[5] ^ bc_6) ^ ad_6) ^ ac_6);
    f_1[6] = (((f_0[6] ^ bc_5) ^ ad_5) ^ ac_5);
    f_1[7] = (((f_0[7] ^ bc_8) ^ ad_8) ^ ac_8);
    f_1[8] = (((f_0[8] ^ bc_7) ^ ad_7) ^ ac_7);
    f_1[9] = (((f_0[9] ^ bc_10) ^ ad_10) ^ ac_10);
    f_1[10] = (((f_0[10] ^ bc_9) ^ ad_9) ^ ac_9);
    f_1[11] = (((f_0[11] ^ bc_12) ^ ad_12) ^ ac_12);
    f_1[12] = (((f_0[12] ^ bc_11) ^ ad_11) ^ ac_11);
  end

  always @(*) begin
    e_2[0] = (((e_1[0] ^ bc_27) ^ ad_27) ^ bd_27);
    e_2[1] = (((e_1[1] ^ bc_26) ^ ad_26) ^ bd_26);
    e_2[2] = (((e_1[2] ^ bc_13) ^ ad_13) ^ bd_13);
    e_2[3] = (((e_1[3] ^ bc_17) ^ ad_17) ^ bd_17);
    e_2[4] = (((e_1[4] ^ bc_16) ^ ad_16) ^ bd_16);
    e_2[5] = (((e_1[5] ^ bc_19) ^ ad_19) ^ bd_19);
    e_2[6] = (((e_1[6] ^ bc_18) ^ ad_18) ^ bd_18);
    e_2[7] = (((e_1[7] ^ bc_21) ^ ad_21) ^ bd_21);
    e_2[8] = (((e_1[8] ^ bc_20) ^ ad_20) ^ bd_20);
    e_2[9] = (((e_1[9] ^ bc_23) ^ ad_23) ^ bd_23);
    e_2[10] = (((e_1[10] ^ bc_22) ^ ad_22) ^ bd_22);
    e_2[11] = (((e_1[11] ^ bc_25) ^ ad_25) ^ bd_25);
    e_2[12] = (((e_1[12] ^ bc_24) ^ ad_24) ^ bd_24);
  end

  always @(*) begin
    f_2[0] = (((f_1[0] ^ bc_27) ^ ad_27) ^ ac_27);
    f_2[1] = (((f_1[1] ^ bc_26) ^ ad_26) ^ ac_26);
    f_2[2] = (((f_1[2] ^ bc_13) ^ ad_13) ^ ac_13);
    f_2[3] = (((f_1[3] ^ bc_17) ^ ad_17) ^ ac_17);
    f_2[4] = (((f_1[4] ^ bc_16) ^ ad_16) ^ ac_16);
    f_2[5] = (((f_1[5] ^ bc_19) ^ ad_19) ^ ac_19);
    f_2[6] = (((f_1[6] ^ bc_18) ^ ad_18) ^ ac_18);
    f_2[7] = (((f_1[7] ^ bc_21) ^ ad_21) ^ ac_21);
    f_2[8] = (((f_1[8] ^ bc_20) ^ ad_20) ^ ac_20);
    f_2[9] = (((f_1[9] ^ bc_23) ^ ad_23) ^ ac_23);
    f_2[10] = (((f_1[10] ^ bc_22) ^ ad_22) ^ ac_22);
    f_2[11] = (((f_1[11] ^ bc_25) ^ ad_25) ^ ac_25);
    f_2[12] = (((f_1[12] ^ bc_24) ^ ad_24) ^ ac_24);
  end

  always @(*) begin
    e_3[0] = (((e_2[0] ^ bc_40) ^ ad_40) ^ bd_40);
    e_3[1] = (((e_2[1] ^ bc_39) ^ ad_39) ^ bd_39);
    e_3[2] = (((e_2[2] ^ bc_43) ^ ad_43) ^ bd_43);
    e_3[3] = (((e_2[3] ^ bc_30) ^ ad_30) ^ bd_30);
    e_3[4] = (((e_2[4] ^ bc_29) ^ ad_29) ^ bd_29);
    e_3[5] = (((e_2[5] ^ bc_32) ^ ad_32) ^ bd_32);
    e_3[6] = (((e_2[6] ^ bc_31) ^ ad_31) ^ bd_31);
    e_3[7] = (((e_2[7] ^ bc_34) ^ ad_34) ^ bd_34);
    e_3[8] = (((e_2[8] ^ bc_33) ^ ad_33) ^ bd_33);
    e_3[9] = (((e_2[9] ^ bc_36) ^ ad_36) ^ bd_36);
    e_3[10] = (((e_2[10] ^ bc_35) ^ ad_35) ^ bd_35);
    e_3[11] = (((e_2[11] ^ bc_38) ^ ad_38) ^ bd_38);
    e_3[12] = (((e_2[12] ^ bc_37) ^ ad_37) ^ bd_37);
  end

  always @(*) begin
    f_3[0] = (((f_2[0] ^ bc_40) ^ ad_40) ^ ac_40);
    f_3[1] = (((f_2[1] ^ bc_39) ^ ad_39) ^ ac_39);
    f_3[2] = (((f_2[2] ^ bc_43) ^ ad_43) ^ ac_43);
    f_3[3] = (((f_2[3] ^ bc_30) ^ ad_30) ^ ac_30);
    f_3[4] = (((f_2[4] ^ bc_29) ^ ad_29) ^ ac_29);
    f_3[5] = (((f_2[5] ^ bc_32) ^ ad_32) ^ ac_32);
    f_3[6] = (((f_2[6] ^ bc_31) ^ ad_31) ^ ac_31);
    f_3[7] = (((f_2[7] ^ bc_34) ^ ad_34) ^ ac_34);
    f_3[8] = (((f_2[8] ^ bc_33) ^ ad_33) ^ ac_33);
    f_3[9] = (((f_2[9] ^ bc_36) ^ ad_36) ^ ac_36);
    f_3[10] = (((f_2[10] ^ bc_35) ^ ad_35) ^ ac_35);
    f_3[11] = (((f_2[11] ^ bc_38) ^ ad_38) ^ ac_38);
    f_3[12] = (((f_2[12] ^ bc_37) ^ ad_37) ^ ac_37);
  end

  always @(*) begin
    e_4[0] = (((e_3[0] ^ bc_53) ^ ad_53) ^ bd_53);
    e_4[1] = (((e_3[1] ^ bc_52) ^ ad_52) ^ bd_52);
    e_4[2] = (((e_3[2] ^ bc_55) ^ ad_55) ^ bd_55);
    e_4[3] = (((e_3[3] ^ bc_54) ^ ad_54) ^ bd_54);
    e_4[4] = (((e_3[4] ^ bc_41) ^ ad_41) ^ bd_41);
    e_4[5] = (((e_3[5] ^ bc_45) ^ ad_45) ^ bd_45);
    e_4[6] = (((e_3[6] ^ bc_44) ^ ad_44) ^ bd_44);
    e_4[7] = (((e_3[7] ^ bc_47) ^ ad_47) ^ bd_47);
    e_4[8] = (((e_3[8] ^ bc_46) ^ ad_46) ^ bd_46);
    e_4[9] = (((e_3[9] ^ bc_49) ^ ad_49) ^ bd_49);
    e_4[10] = (((e_3[10] ^ bc_48) ^ ad_48) ^ bd_48);
    e_4[11] = (((e_3[11] ^ bc_51) ^ ad_51) ^ bd_51);
    e_4[12] = (((e_3[12] ^ bc_50) ^ ad_50) ^ bd_50);
  end

  always @(*) begin
    f_4[0] = (((f_3[0] ^ bc_53) ^ ad_53) ^ ac_53);
    f_4[1] = (((f_3[1] ^ bc_52) ^ ad_52) ^ ac_52);
    f_4[2] = (((f_3[2] ^ bc_55) ^ ad_55) ^ ac_55);
    f_4[3] = (((f_3[3] ^ bc_54) ^ ad_54) ^ ac_54);
    f_4[4] = (((f_3[4] ^ bc_41) ^ ad_41) ^ ac_41);
    f_4[5] = (((f_3[5] ^ bc_45) ^ ad_45) ^ ac_45);
    f_4[6] = (((f_3[6] ^ bc_44) ^ ad_44) ^ ac_44);
    f_4[7] = (((f_3[7] ^ bc_47) ^ ad_47) ^ ac_47);
    f_4[8] = (((f_3[8] ^ bc_46) ^ ad_46) ^ ac_46);
    f_4[9] = (((f_3[9] ^ bc_49) ^ ad_49) ^ ac_49);
    f_4[10] = (((f_3[10] ^ bc_48) ^ ad_48) ^ ac_48);
    f_4[11] = (((f_3[11] ^ bc_51) ^ ad_51) ^ ac_51);
    f_4[12] = (((f_3[12] ^ bc_50) ^ ad_50) ^ ac_50);
  end

  always @(*) begin
    e_5[0] = (((e_4[0] ^ bc_66) ^ ad_66) ^ bd_66);
    e_5[1] = (((e_4[1] ^ bc_65) ^ ad_65) ^ bd_65);
    e_5[2] = (((e_4[2] ^ bc_68) ^ ad_68) ^ bd_68);
    e_5[3] = (((e_4[3] ^ bc_67) ^ ad_67) ^ bd_67);
    e_5[4] = (((e_4[4] ^ bc_71) ^ ad_71) ^ bd_71);
    e_5[5] = (((e_4[5] ^ bc_58) ^ ad_58) ^ bd_58);
    e_5[6] = (((e_4[6] ^ bc_57) ^ ad_57) ^ bd_57);
    e_5[7] = (((e_4[7] ^ bc_60) ^ ad_60) ^ bd_60);
    e_5[8] = (((e_4[8] ^ bc_59) ^ ad_59) ^ bd_59);
    e_5[9] = (((e_4[9] ^ bc_62) ^ ad_62) ^ bd_62);
    e_5[10] = (((e_4[10] ^ bc_61) ^ ad_61) ^ bd_61);
    e_5[11] = (((e_4[11] ^ bc_64) ^ ad_64) ^ bd_64);
    e_5[12] = (((e_4[12] ^ bc_63) ^ ad_63) ^ bd_63);
  end

  always @(*) begin
    f_5[0] = (((f_4[0] ^ bc_66) ^ ad_66) ^ ac_66);
    f_5[1] = (((f_4[1] ^ bc_65) ^ ad_65) ^ ac_65);
    f_5[2] = (((f_4[2] ^ bc_68) ^ ad_68) ^ ac_68);
    f_5[3] = (((f_4[3] ^ bc_67) ^ ad_67) ^ ac_67);
    f_5[4] = (((f_4[4] ^ bc_71) ^ ad_71) ^ ac_71);
    f_5[5] = (((f_4[5] ^ bc_58) ^ ad_58) ^ ac_58);
    f_5[6] = (((f_4[6] ^ bc_57) ^ ad_57) ^ ac_57);
    f_5[7] = (((f_4[7] ^ bc_60) ^ ad_60) ^ ac_60);
    f_5[8] = (((f_4[8] ^ bc_59) ^ ad_59) ^ ac_59);
    f_5[9] = (((f_4[9] ^ bc_62) ^ ad_62) ^ ac_62);
    f_5[10] = (((f_4[10] ^ bc_61) ^ ad_61) ^ ac_61);
    f_5[11] = (((f_4[11] ^ bc_64) ^ ad_64) ^ ac_64);
    f_5[12] = (((f_4[12] ^ bc_63) ^ ad_63) ^ ac_63);
  end

  always @(*) begin
    e_6[0] = (((e_5[0] ^ bc_79) ^ ad_79) ^ bd_79);
    e_6[1] = (((e_5[1] ^ bc_78) ^ ad_78) ^ bd_78);
    e_6[2] = (((e_5[2] ^ bc_81) ^ ad_81) ^ bd_81);
    e_6[3] = (((e_5[3] ^ bc_80) ^ ad_80) ^ bd_80);
    e_6[4] = (((e_5[4] ^ bc_83) ^ ad_83) ^ bd_83);
    e_6[5] = (((e_5[5] ^ bc_82) ^ ad_82) ^ bd_82);
    e_6[6] = (((e_5[6] ^ bc_69) ^ ad_69) ^ bd_69);
    e_6[7] = (((e_5[7] ^ bc_73) ^ ad_73) ^ bd_73);
    e_6[8] = (((e_5[8] ^ bc_72) ^ ad_72) ^ bd_72);
    e_6[9] = (((e_5[9] ^ bc_75) ^ ad_75) ^ bd_75);
    e_6[10] = (((e_5[10] ^ bc_74) ^ ad_74) ^ bd_74);
    e_6[11] = (((e_5[11] ^ bc_77) ^ ad_77) ^ bd_77);
    e_6[12] = (((e_5[12] ^ bc_76) ^ ad_76) ^ bd_76);
  end

  always @(*) begin
    f_6[0] = (((f_5[0] ^ bc_79) ^ ad_79) ^ ac_79);
    f_6[1] = (((f_5[1] ^ bc_78) ^ ad_78) ^ ac_78);
    f_6[2] = (((f_5[2] ^ bc_81) ^ ad_81) ^ ac_81);
    f_6[3] = (((f_5[3] ^ bc_80) ^ ad_80) ^ ac_80);
    f_6[4] = (((f_5[4] ^ bc_83) ^ ad_83) ^ ac_83);
    f_6[5] = (((f_5[5] ^ bc_82) ^ ad_82) ^ ac_82);
    f_6[6] = (((f_5[6] ^ bc_69) ^ ad_69) ^ ac_69);
    f_6[7] = (((f_5[7] ^ bc_73) ^ ad_73) ^ ac_73);
    f_6[8] = (((f_5[8] ^ bc_72) ^ ad_72) ^ ac_72);
    f_6[9] = (((f_5[9] ^ bc_75) ^ ad_75) ^ ac_75);
    f_6[10] = (((f_5[10] ^ bc_74) ^ ad_74) ^ ac_74);
    f_6[11] = (((f_5[11] ^ bc_77) ^ ad_77) ^ ac_77);
    f_6[12] = (((f_5[12] ^ bc_76) ^ ad_76) ^ ac_76);
  end

  always @(*) begin
    e_7[0] = (((e_6[0] ^ bc_92) ^ ad_92) ^ bd_92);
    e_7[1] = (((e_6[1] ^ bc_91) ^ ad_91) ^ bd_91);
    e_7[2] = (((e_6[2] ^ bc_94) ^ ad_94) ^ bd_94);
    e_7[3] = (((e_6[3] ^ bc_93) ^ ad_93) ^ bd_93);
    e_7[4] = (((e_6[4] ^ bc_96) ^ ad_96) ^ bd_96);
    e_7[5] = (((e_6[5] ^ bc_95) ^ ad_95) ^ bd_95);
    e_7[6] = (((e_6[6] ^ bc_99) ^ ad_99) ^ bd_99);
    e_7[7] = (((e_6[7] ^ bc_86) ^ ad_86) ^ bd_86);
    e_7[8] = (((e_6[8] ^ bc_85) ^ ad_85) ^ bd_85);
    e_7[9] = (((e_6[9] ^ bc_88) ^ ad_88) ^ bd_88);
    e_7[10] = (((e_6[10] ^ bc_87) ^ ad_87) ^ bd_87);
    e_7[11] = (((e_6[11] ^ bc_90) ^ ad_90) ^ bd_90);
    e_7[12] = (((e_6[12] ^ bc_89) ^ ad_89) ^ bd_89);
  end

  always @(*) begin
    f_7[0] = (((f_6[0] ^ bc_92) ^ ad_92) ^ ac_92);
    f_7[1] = (((f_6[1] ^ bc_91) ^ ad_91) ^ ac_91);
    f_7[2] = (((f_6[2] ^ bc_94) ^ ad_94) ^ ac_94);
    f_7[3] = (((f_6[3] ^ bc_93) ^ ad_93) ^ ac_93);
    f_7[4] = (((f_6[4] ^ bc_96) ^ ad_96) ^ ac_96);
    f_7[5] = (((f_6[5] ^ bc_95) ^ ad_95) ^ ac_95);
    f_7[6] = (((f_6[6] ^ bc_99) ^ ad_99) ^ ac_99);
    f_7[7] = (((f_6[7] ^ bc_86) ^ ad_86) ^ ac_86);
    f_7[8] = (((f_6[8] ^ bc_85) ^ ad_85) ^ ac_85);
    f_7[9] = (((f_6[9] ^ bc_88) ^ ad_88) ^ ac_88);
    f_7[10] = (((f_6[10] ^ bc_87) ^ ad_87) ^ ac_87);
    f_7[11] = (((f_6[11] ^ bc_90) ^ ad_90) ^ ac_90);
    f_7[12] = (((f_6[12] ^ bc_89) ^ ad_89) ^ ac_89);
  end

  always @(*) begin
    e_8[0] = (((e_7[0] ^ bc_105) ^ ad_105) ^ bd_105);
    e_8[1] = (((e_7[1] ^ bc_104) ^ ad_104) ^ bd_104);
    e_8[2] = (((e_7[2] ^ bc_107) ^ ad_107) ^ bd_107);
    e_8[3] = (((e_7[3] ^ bc_106) ^ ad_106) ^ bd_106);
    e_8[4] = (((e_7[4] ^ bc_109) ^ ad_109) ^ bd_109);
    e_8[5] = (((e_7[5] ^ bc_108) ^ ad_108) ^ bd_108);
    e_8[6] = (((e_7[6] ^ bc_111) ^ ad_111) ^ bd_111);
    e_8[7] = (((e_7[7] ^ bc_110) ^ ad_110) ^ bd_110);
    e_8[8] = (((e_7[8] ^ bc_97) ^ ad_97) ^ bd_97);
    e_8[9] = (((e_7[9] ^ bc_101) ^ ad_101) ^ bd_101);
    e_8[10] = (((e_7[10] ^ bc_100) ^ ad_100) ^ bd_100);
    e_8[11] = (((e_7[11] ^ bc_103) ^ ad_103) ^ bd_103);
    e_8[12] = (((e_7[12] ^ bc_102) ^ ad_102) ^ bd_102);
  end

  always @(*) begin
    f_8[0] = (((f_7[0] ^ bc_105) ^ ad_105) ^ ac_105);
    f_8[1] = (((f_7[1] ^ bc_104) ^ ad_104) ^ ac_104);
    f_8[2] = (((f_7[2] ^ bc_107) ^ ad_107) ^ ac_107);
    f_8[3] = (((f_7[3] ^ bc_106) ^ ad_106) ^ ac_106);
    f_8[4] = (((f_7[4] ^ bc_109) ^ ad_109) ^ ac_109);
    f_8[5] = (((f_7[5] ^ bc_108) ^ ad_108) ^ ac_108);
    f_8[6] = (((f_7[6] ^ bc_111) ^ ad_111) ^ ac_111);
    f_8[7] = (((f_7[7] ^ bc_110) ^ ad_110) ^ ac_110);
    f_8[8] = (((f_7[8] ^ bc_97) ^ ad_97) ^ ac_97);
    f_8[9] = (((f_7[9] ^ bc_101) ^ ad_101) ^ ac_101);
    f_8[10] = (((f_7[10] ^ bc_100) ^ ad_100) ^ ac_100);
    f_8[11] = (((f_7[11] ^ bc_103) ^ ad_103) ^ ac_103);
    f_8[12] = (((f_7[12] ^ bc_102) ^ ad_102) ^ ac_102);
  end

  always @(*) begin
    e_9[0] = (((e_8[0] ^ bc_118) ^ ad_118) ^ bd_118);
    e_9[1] = (((e_8[1] ^ bc_117) ^ ad_117) ^ bd_117);
    e_9[2] = (((e_8[2] ^ bc_120) ^ ad_120) ^ bd_120);
    e_9[3] = (((e_8[3] ^ bc_119) ^ ad_119) ^ bd_119);
    e_9[4] = (((e_8[4] ^ bc_122) ^ ad_122) ^ bd_122);
    e_9[5] = (((e_8[5] ^ bc_121) ^ ad_121) ^ bd_121);
    e_9[6] = (((e_8[6] ^ bc_124) ^ ad_124) ^ bd_124);
    e_9[7] = (((e_8[7] ^ bc_123) ^ ad_123) ^ bd_123);
    e_9[8] = (((e_8[8] ^ bc_127) ^ ad_127) ^ bd_127);
    e_9[9] = (((e_8[9] ^ bc_114) ^ ad_114) ^ bd_114);
    e_9[10] = (((e_8[10] ^ bc_113) ^ ad_113) ^ bd_113);
    e_9[11] = (((e_8[11] ^ bc_116) ^ ad_116) ^ bd_116);
    e_9[12] = (((e_8[12] ^ bc_115) ^ ad_115) ^ bd_115);
  end

  always @(*) begin
    f_9[0] = (((f_8[0] ^ bc_118) ^ ad_118) ^ ac_118);
    f_9[1] = (((f_8[1] ^ bc_117) ^ ad_117) ^ ac_117);
    f_9[2] = (((f_8[2] ^ bc_120) ^ ad_120) ^ ac_120);
    f_9[3] = (((f_8[3] ^ bc_119) ^ ad_119) ^ ac_119);
    f_9[4] = (((f_8[4] ^ bc_122) ^ ad_122) ^ ac_122);
    f_9[5] = (((f_8[5] ^ bc_121) ^ ad_121) ^ ac_121);
    f_9[6] = (((f_8[6] ^ bc_124) ^ ad_124) ^ ac_124);
    f_9[7] = (((f_8[7] ^ bc_123) ^ ad_123) ^ ac_123);
    f_9[8] = (((f_8[8] ^ bc_127) ^ ad_127) ^ ac_127);
    f_9[9] = (((f_8[9] ^ bc_114) ^ ad_114) ^ ac_114);
    f_9[10] = (((f_8[10] ^ bc_113) ^ ad_113) ^ ac_113);
    f_9[11] = (((f_8[11] ^ bc_116) ^ ad_116) ^ ac_116);
    f_9[12] = (((f_8[12] ^ bc_115) ^ ad_115) ^ ac_115);
  end

  always @(*) begin
    e_10[0] = (((e_9[0] ^ bc_131) ^ ad_131) ^ bd_131);
    e_10[1] = (((e_9[1] ^ bc_130) ^ ad_130) ^ bd_130);
    e_10[2] = (((e_9[2] ^ bc_133) ^ ad_133) ^ bd_133);
    e_10[3] = (((e_9[3] ^ bc_132) ^ ad_132) ^ bd_132);
    e_10[4] = (((e_9[4] ^ bc_135) ^ ad_135) ^ bd_135);
    e_10[5] = (((e_9[5] ^ bc_134) ^ ad_134) ^ bd_134);
    e_10[6] = (((e_9[6] ^ bc_137) ^ ad_137) ^ bd_137);
    e_10[7] = (((e_9[7] ^ bc_136) ^ ad_136) ^ bd_136);
    e_10[8] = (((e_9[8] ^ bc_139) ^ ad_139) ^ bd_139);
    e_10[9] = (((e_9[9] ^ bc_138) ^ ad_138) ^ bd_138);
    e_10[10] = (((e_9[10] ^ bc_125) ^ ad_125) ^ bd_125);
    e_10[11] = (((e_9[11] ^ bc_129) ^ ad_129) ^ bd_129);
    e_10[12] = (((e_9[12] ^ bc_128) ^ ad_128) ^ bd_128);
  end

  always @(*) begin
    f_10[0] = (((f_9[0] ^ bc_131) ^ ad_131) ^ ac_131);
    f_10[1] = (((f_9[1] ^ bc_130) ^ ad_130) ^ ac_130);
    f_10[2] = (((f_9[2] ^ bc_133) ^ ad_133) ^ ac_133);
    f_10[3] = (((f_9[3] ^ bc_132) ^ ad_132) ^ ac_132);
    f_10[4] = (((f_9[4] ^ bc_135) ^ ad_135) ^ ac_135);
    f_10[5] = (((f_9[5] ^ bc_134) ^ ad_134) ^ ac_134);
    f_10[6] = (((f_9[6] ^ bc_137) ^ ad_137) ^ ac_137);
    f_10[7] = (((f_9[7] ^ bc_136) ^ ad_136) ^ ac_136);
    f_10[8] = (((f_9[8] ^ bc_139) ^ ad_139) ^ ac_139);
    f_10[9] = (((f_9[9] ^ bc_138) ^ ad_138) ^ ac_138);
    f_10[10] = (((f_9[10] ^ bc_125) ^ ad_125) ^ ac_125);
    f_10[11] = (((f_9[11] ^ bc_129) ^ ad_129) ^ ac_129);
    f_10[12] = (((f_9[12] ^ bc_128) ^ ad_128) ^ ac_128);
  end

  always @(*) begin
    e_11[0] = (((e_10[0] ^ bc_144) ^ ad_144) ^ bd_144);
    e_11[1] = (((e_10[1] ^ bc_143) ^ ad_143) ^ bd_143);
    e_11[2] = (((e_10[2] ^ bc_146) ^ ad_146) ^ bd_146);
    e_11[3] = (((e_10[3] ^ bc_145) ^ ad_145) ^ bd_145);
    e_11[4] = (((e_10[4] ^ bc_148) ^ ad_148) ^ bd_148);
    e_11[5] = (((e_10[5] ^ bc_147) ^ ad_147) ^ bd_147);
    e_11[6] = (((e_10[6] ^ bc_150) ^ ad_150) ^ bd_150);
    e_11[7] = (((e_10[7] ^ bc_149) ^ ad_149) ^ bd_149);
    e_11[8] = (((e_10[8] ^ bc_152) ^ ad_152) ^ bd_152);
    e_11[9] = (((e_10[9] ^ bc_151) ^ ad_151) ^ bd_151);
    e_11[10] = (((e_10[10] ^ bc_155) ^ ad_155) ^ bd_155);
    e_11[11] = (((e_10[11] ^ bc_142) ^ ad_142) ^ bd_142);
    e_11[12] = (((e_10[12] ^ bc_141) ^ ad_141) ^ bd_141);
  end

  always @(*) begin
    f_11[0] = (((f_10[0] ^ bc_144) ^ ad_144) ^ ac_144);
    f_11[1] = (((f_10[1] ^ bc_143) ^ ad_143) ^ ac_143);
    f_11[2] = (((f_10[2] ^ bc_146) ^ ad_146) ^ ac_146);
    f_11[3] = (((f_10[3] ^ bc_145) ^ ad_145) ^ ac_145);
    f_11[4] = (((f_10[4] ^ bc_148) ^ ad_148) ^ ac_148);
    f_11[5] = (((f_10[5] ^ bc_147) ^ ad_147) ^ ac_147);
    f_11[6] = (((f_10[6] ^ bc_150) ^ ad_150) ^ ac_150);
    f_11[7] = (((f_10[7] ^ bc_149) ^ ad_149) ^ ac_149);
    f_11[8] = (((f_10[8] ^ bc_152) ^ ad_152) ^ ac_152);
    f_11[9] = (((f_10[9] ^ bc_151) ^ ad_151) ^ ac_151);
    f_11[10] = (((f_10[10] ^ bc_155) ^ ad_155) ^ ac_155);
    f_11[11] = (((f_10[11] ^ bc_142) ^ ad_142) ^ ac_142);
    f_11[12] = (((f_10[12] ^ bc_141) ^ ad_141) ^ ac_141);
  end

  always @(*) begin
    e_12[0] = (((e_11[0] ^ bc_157) ^ ad_157) ^ bd_157);
    e_12[1] = (((e_11[1] ^ bc_156) ^ ad_156) ^ bd_156);
    e_12[2] = (((e_11[2] ^ bc_159) ^ ad_159) ^ bd_159);
    e_12[3] = (((e_11[3] ^ bc_158) ^ ad_158) ^ bd_158);
    e_12[4] = (((e_11[4] ^ bc_161) ^ ad_161) ^ bd_161);
    e_12[5] = (((e_11[5] ^ bc_160) ^ ad_160) ^ bd_160);
    e_12[6] = (((e_11[6] ^ bc_163) ^ ad_163) ^ bd_163);
    e_12[7] = (((e_11[7] ^ bc_162) ^ ad_162) ^ bd_162);
    e_12[8] = (((e_11[8] ^ bc_165) ^ ad_165) ^ bd_165);
    e_12[9] = (((e_11[9] ^ bc_164) ^ ad_164) ^ bd_164);
    e_12[10] = (((e_11[10] ^ bc_167) ^ ad_167) ^ bd_167);
    e_12[11] = (((e_11[11] ^ bc_166) ^ ad_166) ^ bd_166);
    e_12[12] = (((e_11[12] ^ bc_153) ^ ad_153) ^ bd_153);
  end

  always @(*) begin
    f_12[0] = (((f_11[0] ^ bc_157) ^ ad_157) ^ ac_157);
    f_12[1] = (((f_11[1] ^ bc_156) ^ ad_156) ^ ac_156);
    f_12[2] = (((f_11[2] ^ bc_159) ^ ad_159) ^ ac_159);
    f_12[3] = (((f_11[3] ^ bc_158) ^ ad_158) ^ ac_158);
    f_12[4] = (((f_11[4] ^ bc_161) ^ ad_161) ^ ac_161);
    f_12[5] = (((f_11[5] ^ bc_160) ^ ad_160) ^ ac_160);
    f_12[6] = (((f_11[6] ^ bc_163) ^ ad_163) ^ ac_163);
    f_12[7] = (((f_11[7] ^ bc_162) ^ ad_162) ^ ac_162);
    f_12[8] = (((f_11[8] ^ bc_165) ^ ad_165) ^ ac_165);
    f_12[9] = (((f_11[9] ^ bc_164) ^ ad_164) ^ ac_164);
    f_12[10] = (((f_11[10] ^ bc_167) ^ ad_167) ^ ac_167);
    f_12[11] = (((f_11[11] ^ bc_166) ^ ad_166) ^ ac_166);
    f_12[12] = (((f_11[12] ^ bc_153) ^ ad_153) ^ ac_153);
  end

  assign io_z_0 = {e_12[0],f_12[0]};
  assign io_z_1 = {e_12[1],f_12[1]};
  assign io_z_2 = {e_12[2],f_12[2]};
  assign io_z_3 = {e_12[3],f_12[3]};
  assign io_z_4 = {e_12[4],f_12[4]};
  assign io_z_5 = {e_12[5],f_12[5]};
  assign io_z_6 = {e_12[6],f_12[6]};
  assign io_z_7 = {e_12[7],f_12[7]};
  assign io_z_8 = {e_12[8],f_12[8]};
  assign io_z_9 = {e_12[9],f_12[9]};
  assign io_z_10 = {e_12[10],f_12[10]};
  assign io_z_11 = {e_12[11],f_12[11]};
  assign io_z_12 = {e_12[12],f_12[12]};

endmodule
