-- Generator : SpinalHDL v1.6.2    git head : 685405804ac0fa51f884fe0ee6813ba6f1f31e4e
-- Component : aesEncrypt_Unrolled
-- Git hash  : 685405804ac0fa51f884fe0ee6813ba6f1f31e4e

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;

package pkg_enum is

end pkg_enum;

library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

package pkg_scala2hdl is
  function pkg_extract (that : std_logic_vector; bitId : integer) return std_logic;
  function pkg_extract (that : std_logic_vector; base : unsigned; size : integer) return std_logic_vector;
  function pkg_cat (a : std_logic_vector; b : std_logic_vector) return std_logic_vector;
  function pkg_not (value : std_logic_vector) return std_logic_vector;
  function pkg_extract (that : unsigned; bitId : integer) return std_logic;
  function pkg_extract (that : unsigned; base : unsigned; size : integer) return unsigned;
  function pkg_cat (a : unsigned; b : unsigned) return unsigned;
  function pkg_not (value : unsigned) return unsigned;
  function pkg_extract (that : signed; bitId : integer) return std_logic;
  function pkg_extract (that : signed; base : unsigned; size : integer) return signed;
  function pkg_cat (a : signed; b : signed) return signed;
  function pkg_not (value : signed) return signed;

  function pkg_mux (sel : std_logic; one : std_logic; zero : std_logic) return std_logic;
  function pkg_mux (sel : std_logic; one : std_logic_vector; zero : std_logic_vector) return std_logic_vector;
  function pkg_mux (sel : std_logic; one : unsigned; zero : unsigned) return unsigned;
  function pkg_mux (sel : std_logic; one : signed; zero : signed) return signed;

  function pkg_toStdLogic (value : boolean) return std_logic;
  function pkg_toStdLogicVector (value : std_logic) return std_logic_vector;
  function pkg_toUnsigned (value : std_logic) return unsigned;
  function pkg_toSigned (value : std_logic) return signed;
  function pkg_stdLogicVector (lit : std_logic_vector) return std_logic_vector;
  function pkg_unsigned (lit : unsigned) return unsigned;
  function pkg_signed (lit : signed) return signed;

  function pkg_resize (that : std_logic_vector; width : integer) return std_logic_vector;
  function pkg_resize (that : unsigned; width : integer) return unsigned;
  function pkg_resize (that : signed; width : integer) return signed;

  function pkg_extract (that : std_logic_vector; high : integer; low : integer) return std_logic_vector;
  function pkg_extract (that : unsigned; high : integer; low : integer) return unsigned;
  function pkg_extract (that : signed; high : integer; low : integer) return signed;

  function pkg_shiftRight (that : std_logic_vector; size : natural) return std_logic_vector;
  function pkg_shiftRight (that : std_logic_vector; size : unsigned) return std_logic_vector;
  function pkg_shiftLeft (that : std_logic_vector; size : natural) return std_logic_vector;
  function pkg_shiftLeft (that : std_logic_vector; size : unsigned) return std_logic_vector;

  function pkg_shiftRight (that : unsigned; size : natural) return unsigned;
  function pkg_shiftRight (that : unsigned; size : unsigned) return unsigned;
  function pkg_shiftLeft (that : unsigned; size : natural) return unsigned;
  function pkg_shiftLeft (that : unsigned; size : unsigned) return unsigned;

  function pkg_shiftRight (that : signed; size : natural) return signed;
  function pkg_shiftRight (that : signed; size : unsigned) return signed;
  function pkg_shiftLeft (that : signed; size : natural) return signed;
  function pkg_shiftLeft (that : signed; size : unsigned; w : integer) return signed;

  function pkg_rotateLeft (that : std_logic_vector; size : unsigned) return std_logic_vector;
end  pkg_scala2hdl;

package body pkg_scala2hdl is
  function pkg_extract (that : std_logic_vector; bitId : integer) return std_logic is
    alias temp : std_logic_vector(that'length-1 downto 0) is that;
  begin
    return temp(bitId);
  end pkg_extract;

  function pkg_extract (that : std_logic_vector; base : unsigned; size : integer) return std_logic_vector is
    alias temp : std_logic_vector(that'length-1 downto 0) is that;    constant elementCount : integer := temp'length - size + 1;
    type tableType is array (0 to elementCount-1) of std_logic_vector(size-1 downto 0);
    variable table : tableType;
  begin
    for i in 0 to elementCount-1 loop
      table(i) := temp(i + size - 1 downto i);
    end loop;
    return table(to_integer(base));
  end pkg_extract;

  function pkg_cat (a : std_logic_vector; b : std_logic_vector) return std_logic_vector is
    variable cat : std_logic_vector(a'length + b'length-1 downto 0);
  begin
    cat := a & b;
    return cat;
  end pkg_cat;

  function pkg_not (value : std_logic_vector) return std_logic_vector is
    variable ret : std_logic_vector(value'length-1 downto 0);
  begin
    ret := not value;
    return ret;
  end pkg_not;

  function pkg_extract (that : unsigned; bitId : integer) return std_logic is
    alias temp : unsigned(that'length-1 downto 0) is that;
  begin
    return temp(bitId);
  end pkg_extract;

  function pkg_extract (that : unsigned; base : unsigned; size : integer) return unsigned is
    alias temp : unsigned(that'length-1 downto 0) is that;    constant elementCount : integer := temp'length - size + 1;
    type tableType is array (0 to elementCount-1) of unsigned(size-1 downto 0);
    variable table : tableType;
  begin
    for i in 0 to elementCount-1 loop
      table(i) := temp(i + size - 1 downto i);
    end loop;
    return table(to_integer(base));
  end pkg_extract;

  function pkg_cat (a : unsigned; b : unsigned) return unsigned is
    variable cat : unsigned(a'length + b'length-1 downto 0);
  begin
    cat := a & b;
    return cat;
  end pkg_cat;

  function pkg_not (value : unsigned) return unsigned is
    variable ret : unsigned(value'length-1 downto 0);
  begin
    ret := not value;
    return ret;
  end pkg_not;

  function pkg_extract (that : signed; bitId : integer) return std_logic is
    alias temp : signed(that'length-1 downto 0) is that;
  begin
    return temp(bitId);
  end pkg_extract;

  function pkg_extract (that : signed; base : unsigned; size : integer) return signed is
    alias temp : signed(that'length-1 downto 0) is that;    constant elementCount : integer := temp'length - size + 1;
    type tableType is array (0 to elementCount-1) of signed(size-1 downto 0);
    variable table : tableType;
  begin
    for i in 0 to elementCount-1 loop
      table(i) := temp(i + size - 1 downto i);
    end loop;
    return table(to_integer(base));
  end pkg_extract;

  function pkg_cat (a : signed; b : signed) return signed is
    variable cat : signed(a'length + b'length-1 downto 0);
  begin
    cat := a & b;
    return cat;
  end pkg_cat;

  function pkg_not (value : signed) return signed is
    variable ret : signed(value'length-1 downto 0);
  begin
    ret := not value;
    return ret;
  end pkg_not;


  -- unsigned shifts
  function pkg_shiftRight (that : unsigned; size : natural) return unsigned is
    variable ret : unsigned(that'length-1 downto 0);
  begin
    if size >= that'length then
      return "";
    else
      ret := shift_right(that,size);
      return ret(that'length-1-size downto 0);
    end if;
  end pkg_shiftRight;

  function pkg_shiftRight (that : unsigned; size : unsigned) return unsigned is
    variable ret : unsigned(that'length-1 downto 0);
  begin
    ret := shift_right(that,to_integer(size));
    return ret;
  end pkg_shiftRight;

  function pkg_shiftLeft (that : unsigned; size : natural) return unsigned is
  begin
    return shift_left(resize(that,that'length + size),size);
  end pkg_shiftLeft;

  function pkg_shiftLeft (that : unsigned; size : unsigned) return unsigned is
  begin
    return shift_left(resize(that,that'length + 2**size'length - 1),to_integer(size));
  end pkg_shiftLeft;

  -- std_logic_vector shifts
  function pkg_shiftRight (that : std_logic_vector; size : natural) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftRight(unsigned(that),size));
  end pkg_shiftRight;

  function pkg_shiftRight (that : std_logic_vector; size : unsigned) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftRight(unsigned(that),size));
  end pkg_shiftRight;

  function pkg_shiftLeft (that : std_logic_vector; size : natural) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftLeft(unsigned(that),size));
  end pkg_shiftLeft;

  function pkg_shiftLeft (that : std_logic_vector; size : unsigned) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftLeft(unsigned(that),size));
  end pkg_shiftLeft;

  -- signed shifts
  function pkg_shiftRight (that : signed; size : natural) return signed is
  begin
    return signed(pkg_shiftRight(unsigned(that),size));
  end pkg_shiftRight;

  function pkg_shiftRight (that : signed; size : unsigned) return signed is
  begin
    return shift_right(that,to_integer(size));
  end pkg_shiftRight;

  function pkg_shiftLeft (that : signed; size : natural) return signed is
  begin
    return signed(pkg_shiftLeft(unsigned(that),size));
  end pkg_shiftLeft;

  function pkg_shiftLeft (that : signed; size : unsigned; w : integer) return signed is
  begin
    return shift_left(resize(that,w),to_integer(size));
  end pkg_shiftLeft;

  function pkg_rotateLeft (that : std_logic_vector; size : unsigned) return std_logic_vector is
  begin
    return std_logic_vector(rotate_left(unsigned(that),to_integer(size)));
  end pkg_rotateLeft;

  function pkg_extract (that : std_logic_vector; high : integer; low : integer) return std_logic_vector is
    alias temp : std_logic_vector(that'length-1 downto 0) is that;
  begin
    return temp(high downto low);
  end pkg_extract;

  function pkg_extract (that : unsigned; high : integer; low : integer) return unsigned is
    alias temp : unsigned(that'length-1 downto 0) is that;
  begin
    return temp(high downto low);
  end pkg_extract;

  function pkg_extract (that : signed; high : integer; low : integer) return signed is
    alias temp : signed(that'length-1 downto 0) is that;
  begin
    return temp(high downto low);
  end pkg_extract;

  function pkg_mux (sel : std_logic; one : std_logic; zero : std_logic) return std_logic is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : std_logic_vector; zero : std_logic_vector) return std_logic_vector is
    variable ret : std_logic_vector(zero'range);
  begin
    if sel = '1' then
      ret := one;
    else
      ret := zero;
    end if;
    return ret;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : unsigned; zero : unsigned) return unsigned is
    variable ret : unsigned(zero'range);
  begin
    if sel = '1' then
      ret := one;
    else
      ret := zero;
    end if;
    return ret;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : signed; zero : signed) return signed is
    variable ret : signed(zero'range);
  begin
    if sel = '1' then
      ret := one;
    else
      ret := zero;
    end if;
    return ret;
  end pkg_mux;

  function pkg_toStdLogic (value : boolean) return std_logic is
  begin
    if value = true then
      return '1';
    else
      return '0';
    end if;
  end pkg_toStdLogic;

  function pkg_toStdLogicVector (value : std_logic) return std_logic_vector is
    variable ret : std_logic_vector(0 downto 0);
  begin
    ret(0) := value;
    return ret;
  end pkg_toStdLogicVector;

  function pkg_toUnsigned (value : std_logic) return unsigned is
    variable ret : unsigned(0 downto 0);
  begin
    ret(0) := value;
    return ret;
  end pkg_toUnsigned;

  function pkg_toSigned (value : std_logic) return signed is
    variable ret : signed(0 downto 0);
  begin
    ret(0) := value;
    return ret;
  end pkg_toSigned;

  function pkg_stdLogicVector (lit : std_logic_vector) return std_logic_vector is
    alias ret : std_logic_vector(lit'length-1 downto 0) is lit;
  begin
    return ret;
  end pkg_stdLogicVector;

  function pkg_unsigned (lit : unsigned) return unsigned is
    alias ret : unsigned(lit'length-1 downto 0) is lit;
  begin
    return ret;
  end pkg_unsigned;

  function pkg_signed (lit : signed) return signed is
    alias ret : signed(lit'length-1 downto 0) is lit;
  begin
    return ret;
  end pkg_signed;

  function pkg_resize (that : std_logic_vector; width : integer) return std_logic_vector is
  begin
    return std_logic_vector(resize(unsigned(that),width));
  end pkg_resize;

  function pkg_resize (that : unsigned; width : integer) return unsigned is
    variable ret : unsigned(width-1 downto 0);
  begin
    if that'length = 0 then
       ret := (others => '0');
    else
       ret := resize(that,width);
    end if;
    return ret;
  end pkg_resize;
  function pkg_resize (that : signed; width : integer) return signed is
    alias temp : signed(that'length-1 downto 0) is that;
    variable ret : signed(width-1 downto 0);
  begin
    if temp'length = 0 then
       ret := (others => '0');
    elsif temp'length >= width then
       ret := temp(width-1 downto 0);
    else
       ret := resize(temp,width);
    end if;
    return ret;
  end pkg_resize;
end pkg_scala2hdl;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity SubByte is
  port(
    io_b : in std_logic_vector(7 downto 0);
    io_ret : out std_logic_vector(7 downto 0)
  );
end SubByte;

architecture arch of SubByte is

  signal zz_io_ret : std_logic_vector(7 downto 0);
begin
  process(io_b)
  begin
    case io_b is
      when "00000000" =>
        zz_io_ret <= pkg_stdLogicVector("01100011");
      when "00000001" =>
        zz_io_ret <= pkg_stdLogicVector("01111100");
      when "00000010" =>
        zz_io_ret <= pkg_stdLogicVector("01110111");
      when "00000011" =>
        zz_io_ret <= pkg_stdLogicVector("01111011");
      when "00000100" =>
        zz_io_ret <= pkg_stdLogicVector("11110010");
      when "00000101" =>
        zz_io_ret <= pkg_stdLogicVector("01101011");
      when "00000110" =>
        zz_io_ret <= pkg_stdLogicVector("01101111");
      when "00000111" =>
        zz_io_ret <= pkg_stdLogicVector("11000101");
      when "00001000" =>
        zz_io_ret <= pkg_stdLogicVector("00110000");
      when "00001001" =>
        zz_io_ret <= pkg_stdLogicVector("00000001");
      when "00001010" =>
        zz_io_ret <= pkg_stdLogicVector("01100111");
      when "00001011" =>
        zz_io_ret <= pkg_stdLogicVector("00101011");
      when "00001100" =>
        zz_io_ret <= pkg_stdLogicVector("11111110");
      when "00001101" =>
        zz_io_ret <= pkg_stdLogicVector("11010111");
      when "00001110" =>
        zz_io_ret <= pkg_stdLogicVector("10101011");
      when "00001111" =>
        zz_io_ret <= pkg_stdLogicVector("01110110");
      when "00010000" =>
        zz_io_ret <= pkg_stdLogicVector("11001010");
      when "00010001" =>
        zz_io_ret <= pkg_stdLogicVector("10000010");
      when "00010010" =>
        zz_io_ret <= pkg_stdLogicVector("11001001");
      when "00010011" =>
        zz_io_ret <= pkg_stdLogicVector("01111101");
      when "00010100" =>
        zz_io_ret <= pkg_stdLogicVector("11111010");
      when "00010101" =>
        zz_io_ret <= pkg_stdLogicVector("01011001");
      when "00010110" =>
        zz_io_ret <= pkg_stdLogicVector("01000111");
      when "00010111" =>
        zz_io_ret <= pkg_stdLogicVector("11110000");
      when "00011000" =>
        zz_io_ret <= pkg_stdLogicVector("10101101");
      when "00011001" =>
        zz_io_ret <= pkg_stdLogicVector("11010100");
      when "00011010" =>
        zz_io_ret <= pkg_stdLogicVector("10100010");
      when "00011011" =>
        zz_io_ret <= pkg_stdLogicVector("10101111");
      when "00011100" =>
        zz_io_ret <= pkg_stdLogicVector("10011100");
      when "00011101" =>
        zz_io_ret <= pkg_stdLogicVector("10100100");
      when "00011110" =>
        zz_io_ret <= pkg_stdLogicVector("01110010");
      when "00011111" =>
        zz_io_ret <= pkg_stdLogicVector("11000000");
      when "00100000" =>
        zz_io_ret <= pkg_stdLogicVector("10110111");
      when "00100001" =>
        zz_io_ret <= pkg_stdLogicVector("11111101");
      when "00100010" =>
        zz_io_ret <= pkg_stdLogicVector("10010011");
      when "00100011" =>
        zz_io_ret <= pkg_stdLogicVector("00100110");
      when "00100100" =>
        zz_io_ret <= pkg_stdLogicVector("00110110");
      when "00100101" =>
        zz_io_ret <= pkg_stdLogicVector("00111111");
      when "00100110" =>
        zz_io_ret <= pkg_stdLogicVector("11110111");
      when "00100111" =>
        zz_io_ret <= pkg_stdLogicVector("11001100");
      when "00101000" =>
        zz_io_ret <= pkg_stdLogicVector("00110100");
      when "00101001" =>
        zz_io_ret <= pkg_stdLogicVector("10100101");
      when "00101010" =>
        zz_io_ret <= pkg_stdLogicVector("11100101");
      when "00101011" =>
        zz_io_ret <= pkg_stdLogicVector("11110001");
      when "00101100" =>
        zz_io_ret <= pkg_stdLogicVector("01110001");
      when "00101101" =>
        zz_io_ret <= pkg_stdLogicVector("11011000");
      when "00101110" =>
        zz_io_ret <= pkg_stdLogicVector("00110001");
      when "00101111" =>
        zz_io_ret <= pkg_stdLogicVector("00010101");
      when "00110000" =>
        zz_io_ret <= pkg_stdLogicVector("00000100");
      when "00110001" =>
        zz_io_ret <= pkg_stdLogicVector("11000111");
      when "00110010" =>
        zz_io_ret <= pkg_stdLogicVector("00100011");
      when "00110011" =>
        zz_io_ret <= pkg_stdLogicVector("11000011");
      when "00110100" =>
        zz_io_ret <= pkg_stdLogicVector("00011000");
      when "00110101" =>
        zz_io_ret <= pkg_stdLogicVector("10010110");
      when "00110110" =>
        zz_io_ret <= pkg_stdLogicVector("00000101");
      when "00110111" =>
        zz_io_ret <= pkg_stdLogicVector("10011010");
      when "00111000" =>
        zz_io_ret <= pkg_stdLogicVector("00000111");
      when "00111001" =>
        zz_io_ret <= pkg_stdLogicVector("00010010");
      when "00111010" =>
        zz_io_ret <= pkg_stdLogicVector("10000000");
      when "00111011" =>
        zz_io_ret <= pkg_stdLogicVector("11100010");
      when "00111100" =>
        zz_io_ret <= pkg_stdLogicVector("11101011");
      when "00111101" =>
        zz_io_ret <= pkg_stdLogicVector("00100111");
      when "00111110" =>
        zz_io_ret <= pkg_stdLogicVector("10110010");
      when "00111111" =>
        zz_io_ret <= pkg_stdLogicVector("01110101");
      when "01000000" =>
        zz_io_ret <= pkg_stdLogicVector("00001001");
      when "01000001" =>
        zz_io_ret <= pkg_stdLogicVector("10000011");
      when "01000010" =>
        zz_io_ret <= pkg_stdLogicVector("00101100");
      when "01000011" =>
        zz_io_ret <= pkg_stdLogicVector("00011010");
      when "01000100" =>
        zz_io_ret <= pkg_stdLogicVector("00011011");
      when "01000101" =>
        zz_io_ret <= pkg_stdLogicVector("01101110");
      when "01000110" =>
        zz_io_ret <= pkg_stdLogicVector("01011010");
      when "01000111" =>
        zz_io_ret <= pkg_stdLogicVector("10100000");
      when "01001000" =>
        zz_io_ret <= pkg_stdLogicVector("01010010");
      when "01001001" =>
        zz_io_ret <= pkg_stdLogicVector("00111011");
      when "01001010" =>
        zz_io_ret <= pkg_stdLogicVector("11010110");
      when "01001011" =>
        zz_io_ret <= pkg_stdLogicVector("10110011");
      when "01001100" =>
        zz_io_ret <= pkg_stdLogicVector("00101001");
      when "01001101" =>
        zz_io_ret <= pkg_stdLogicVector("11100011");
      when "01001110" =>
        zz_io_ret <= pkg_stdLogicVector("00101111");
      when "01001111" =>
        zz_io_ret <= pkg_stdLogicVector("10000100");
      when "01010000" =>
        zz_io_ret <= pkg_stdLogicVector("01010011");
      when "01010001" =>
        zz_io_ret <= pkg_stdLogicVector("11010001");
      when "01010010" =>
        zz_io_ret <= pkg_stdLogicVector("00000000");
      when "01010011" =>
        zz_io_ret <= pkg_stdLogicVector("11101101");
      when "01010100" =>
        zz_io_ret <= pkg_stdLogicVector("00100000");
      when "01010101" =>
        zz_io_ret <= pkg_stdLogicVector("11111100");
      when "01010110" =>
        zz_io_ret <= pkg_stdLogicVector("10110001");
      when "01010111" =>
        zz_io_ret <= pkg_stdLogicVector("01011011");
      when "01011000" =>
        zz_io_ret <= pkg_stdLogicVector("01101010");
      when "01011001" =>
        zz_io_ret <= pkg_stdLogicVector("11001011");
      when "01011010" =>
        zz_io_ret <= pkg_stdLogicVector("10111110");
      when "01011011" =>
        zz_io_ret <= pkg_stdLogicVector("00111001");
      when "01011100" =>
        zz_io_ret <= pkg_stdLogicVector("01001010");
      when "01011101" =>
        zz_io_ret <= pkg_stdLogicVector("01001100");
      when "01011110" =>
        zz_io_ret <= pkg_stdLogicVector("01011000");
      when "01011111" =>
        zz_io_ret <= pkg_stdLogicVector("11001111");
      when "01100000" =>
        zz_io_ret <= pkg_stdLogicVector("11010000");
      when "01100001" =>
        zz_io_ret <= pkg_stdLogicVector("11101111");
      when "01100010" =>
        zz_io_ret <= pkg_stdLogicVector("10101010");
      when "01100011" =>
        zz_io_ret <= pkg_stdLogicVector("11111011");
      when "01100100" =>
        zz_io_ret <= pkg_stdLogicVector("01000011");
      when "01100101" =>
        zz_io_ret <= pkg_stdLogicVector("01001101");
      when "01100110" =>
        zz_io_ret <= pkg_stdLogicVector("00110011");
      when "01100111" =>
        zz_io_ret <= pkg_stdLogicVector("10000101");
      when "01101000" =>
        zz_io_ret <= pkg_stdLogicVector("01000101");
      when "01101001" =>
        zz_io_ret <= pkg_stdLogicVector("11111001");
      when "01101010" =>
        zz_io_ret <= pkg_stdLogicVector("00000010");
      when "01101011" =>
        zz_io_ret <= pkg_stdLogicVector("01111111");
      when "01101100" =>
        zz_io_ret <= pkg_stdLogicVector("01010000");
      when "01101101" =>
        zz_io_ret <= pkg_stdLogicVector("00111100");
      when "01101110" =>
        zz_io_ret <= pkg_stdLogicVector("10011111");
      when "01101111" =>
        zz_io_ret <= pkg_stdLogicVector("10101000");
      when "01110000" =>
        zz_io_ret <= pkg_stdLogicVector("01010001");
      when "01110001" =>
        zz_io_ret <= pkg_stdLogicVector("10100011");
      when "01110010" =>
        zz_io_ret <= pkg_stdLogicVector("01000000");
      when "01110011" =>
        zz_io_ret <= pkg_stdLogicVector("10001111");
      when "01110100" =>
        zz_io_ret <= pkg_stdLogicVector("10010010");
      when "01110101" =>
        zz_io_ret <= pkg_stdLogicVector("10011101");
      when "01110110" =>
        zz_io_ret <= pkg_stdLogicVector("00111000");
      when "01110111" =>
        zz_io_ret <= pkg_stdLogicVector("11110101");
      when "01111000" =>
        zz_io_ret <= pkg_stdLogicVector("10111100");
      when "01111001" =>
        zz_io_ret <= pkg_stdLogicVector("10110110");
      when "01111010" =>
        zz_io_ret <= pkg_stdLogicVector("11011010");
      when "01111011" =>
        zz_io_ret <= pkg_stdLogicVector("00100001");
      when "01111100" =>
        zz_io_ret <= pkg_stdLogicVector("00010000");
      when "01111101" =>
        zz_io_ret <= pkg_stdLogicVector("11111111");
      when "01111110" =>
        zz_io_ret <= pkg_stdLogicVector("11110011");
      when "01111111" =>
        zz_io_ret <= pkg_stdLogicVector("11010010");
      when "10000000" =>
        zz_io_ret <= pkg_stdLogicVector("11001101");
      when "10000001" =>
        zz_io_ret <= pkg_stdLogicVector("00001100");
      when "10000010" =>
        zz_io_ret <= pkg_stdLogicVector("00010011");
      when "10000011" =>
        zz_io_ret <= pkg_stdLogicVector("11101100");
      when "10000100" =>
        zz_io_ret <= pkg_stdLogicVector("01011111");
      when "10000101" =>
        zz_io_ret <= pkg_stdLogicVector("10010111");
      when "10000110" =>
        zz_io_ret <= pkg_stdLogicVector("01000100");
      when "10000111" =>
        zz_io_ret <= pkg_stdLogicVector("00010111");
      when "10001000" =>
        zz_io_ret <= pkg_stdLogicVector("11000100");
      when "10001001" =>
        zz_io_ret <= pkg_stdLogicVector("10100111");
      when "10001010" =>
        zz_io_ret <= pkg_stdLogicVector("01111110");
      when "10001011" =>
        zz_io_ret <= pkg_stdLogicVector("00111101");
      when "10001100" =>
        zz_io_ret <= pkg_stdLogicVector("01100100");
      when "10001101" =>
        zz_io_ret <= pkg_stdLogicVector("01011101");
      when "10001110" =>
        zz_io_ret <= pkg_stdLogicVector("00011001");
      when "10001111" =>
        zz_io_ret <= pkg_stdLogicVector("01110011");
      when "10010000" =>
        zz_io_ret <= pkg_stdLogicVector("01100000");
      when "10010001" =>
        zz_io_ret <= pkg_stdLogicVector("10000001");
      when "10010010" =>
        zz_io_ret <= pkg_stdLogicVector("01001111");
      when "10010011" =>
        zz_io_ret <= pkg_stdLogicVector("11011100");
      when "10010100" =>
        zz_io_ret <= pkg_stdLogicVector("00100010");
      when "10010101" =>
        zz_io_ret <= pkg_stdLogicVector("00101010");
      when "10010110" =>
        zz_io_ret <= pkg_stdLogicVector("10010000");
      when "10010111" =>
        zz_io_ret <= pkg_stdLogicVector("10001000");
      when "10011000" =>
        zz_io_ret <= pkg_stdLogicVector("01000110");
      when "10011001" =>
        zz_io_ret <= pkg_stdLogicVector("11101110");
      when "10011010" =>
        zz_io_ret <= pkg_stdLogicVector("10111000");
      when "10011011" =>
        zz_io_ret <= pkg_stdLogicVector("00010100");
      when "10011100" =>
        zz_io_ret <= pkg_stdLogicVector("11011110");
      when "10011101" =>
        zz_io_ret <= pkg_stdLogicVector("01011110");
      when "10011110" =>
        zz_io_ret <= pkg_stdLogicVector("00001011");
      when "10011111" =>
        zz_io_ret <= pkg_stdLogicVector("11011011");
      when "10100000" =>
        zz_io_ret <= pkg_stdLogicVector("11100000");
      when "10100001" =>
        zz_io_ret <= pkg_stdLogicVector("00110010");
      when "10100010" =>
        zz_io_ret <= pkg_stdLogicVector("00111010");
      when "10100011" =>
        zz_io_ret <= pkg_stdLogicVector("00001010");
      when "10100100" =>
        zz_io_ret <= pkg_stdLogicVector("01001001");
      when "10100101" =>
        zz_io_ret <= pkg_stdLogicVector("00000110");
      when "10100110" =>
        zz_io_ret <= pkg_stdLogicVector("00100100");
      when "10100111" =>
        zz_io_ret <= pkg_stdLogicVector("01011100");
      when "10101000" =>
        zz_io_ret <= pkg_stdLogicVector("11000010");
      when "10101001" =>
        zz_io_ret <= pkg_stdLogicVector("11010011");
      when "10101010" =>
        zz_io_ret <= pkg_stdLogicVector("10101100");
      when "10101011" =>
        zz_io_ret <= pkg_stdLogicVector("01100010");
      when "10101100" =>
        zz_io_ret <= pkg_stdLogicVector("10010001");
      when "10101101" =>
        zz_io_ret <= pkg_stdLogicVector("10010101");
      when "10101110" =>
        zz_io_ret <= pkg_stdLogicVector("11100100");
      when "10101111" =>
        zz_io_ret <= pkg_stdLogicVector("01111001");
      when "10110000" =>
        zz_io_ret <= pkg_stdLogicVector("11100111");
      when "10110001" =>
        zz_io_ret <= pkg_stdLogicVector("11001000");
      when "10110010" =>
        zz_io_ret <= pkg_stdLogicVector("00110111");
      when "10110011" =>
        zz_io_ret <= pkg_stdLogicVector("01101101");
      when "10110100" =>
        zz_io_ret <= pkg_stdLogicVector("10001101");
      when "10110101" =>
        zz_io_ret <= pkg_stdLogicVector("11010101");
      when "10110110" =>
        zz_io_ret <= pkg_stdLogicVector("01001110");
      when "10110111" =>
        zz_io_ret <= pkg_stdLogicVector("10101001");
      when "10111000" =>
        zz_io_ret <= pkg_stdLogicVector("01101100");
      when "10111001" =>
        zz_io_ret <= pkg_stdLogicVector("01010110");
      when "10111010" =>
        zz_io_ret <= pkg_stdLogicVector("11110100");
      when "10111011" =>
        zz_io_ret <= pkg_stdLogicVector("11101010");
      when "10111100" =>
        zz_io_ret <= pkg_stdLogicVector("01100101");
      when "10111101" =>
        zz_io_ret <= pkg_stdLogicVector("01111010");
      when "10111110" =>
        zz_io_ret <= pkg_stdLogicVector("10101110");
      when "10111111" =>
        zz_io_ret <= pkg_stdLogicVector("00001000");
      when "11000000" =>
        zz_io_ret <= pkg_stdLogicVector("10111010");
      when "11000001" =>
        zz_io_ret <= pkg_stdLogicVector("01111000");
      when "11000010" =>
        zz_io_ret <= pkg_stdLogicVector("00100101");
      when "11000011" =>
        zz_io_ret <= pkg_stdLogicVector("00101110");
      when "11000100" =>
        zz_io_ret <= pkg_stdLogicVector("00011100");
      when "11000101" =>
        zz_io_ret <= pkg_stdLogicVector("10100110");
      when "11000110" =>
        zz_io_ret <= pkg_stdLogicVector("10110100");
      when "11000111" =>
        zz_io_ret <= pkg_stdLogicVector("11000110");
      when "11001000" =>
        zz_io_ret <= pkg_stdLogicVector("11101000");
      when "11001001" =>
        zz_io_ret <= pkg_stdLogicVector("11011101");
      when "11001010" =>
        zz_io_ret <= pkg_stdLogicVector("01110100");
      when "11001011" =>
        zz_io_ret <= pkg_stdLogicVector("00011111");
      when "11001100" =>
        zz_io_ret <= pkg_stdLogicVector("01001011");
      when "11001101" =>
        zz_io_ret <= pkg_stdLogicVector("10111101");
      when "11001110" =>
        zz_io_ret <= pkg_stdLogicVector("10001011");
      when "11001111" =>
        zz_io_ret <= pkg_stdLogicVector("10001010");
      when "11010000" =>
        zz_io_ret <= pkg_stdLogicVector("01110000");
      when "11010001" =>
        zz_io_ret <= pkg_stdLogicVector("00111110");
      when "11010010" =>
        zz_io_ret <= pkg_stdLogicVector("10110101");
      when "11010011" =>
        zz_io_ret <= pkg_stdLogicVector("01100110");
      when "11010100" =>
        zz_io_ret <= pkg_stdLogicVector("01001000");
      when "11010101" =>
        zz_io_ret <= pkg_stdLogicVector("00000011");
      when "11010110" =>
        zz_io_ret <= pkg_stdLogicVector("11110110");
      when "11010111" =>
        zz_io_ret <= pkg_stdLogicVector("00001110");
      when "11011000" =>
        zz_io_ret <= pkg_stdLogicVector("01100001");
      when "11011001" =>
        zz_io_ret <= pkg_stdLogicVector("00110101");
      when "11011010" =>
        zz_io_ret <= pkg_stdLogicVector("01010111");
      when "11011011" =>
        zz_io_ret <= pkg_stdLogicVector("10111001");
      when "11011100" =>
        zz_io_ret <= pkg_stdLogicVector("10000110");
      when "11011101" =>
        zz_io_ret <= pkg_stdLogicVector("11000001");
      when "11011110" =>
        zz_io_ret <= pkg_stdLogicVector("00011101");
      when "11011111" =>
        zz_io_ret <= pkg_stdLogicVector("10011110");
      when "11100000" =>
        zz_io_ret <= pkg_stdLogicVector("11100001");
      when "11100001" =>
        zz_io_ret <= pkg_stdLogicVector("11111000");
      when "11100010" =>
        zz_io_ret <= pkg_stdLogicVector("10011000");
      when "11100011" =>
        zz_io_ret <= pkg_stdLogicVector("00010001");
      when "11100100" =>
        zz_io_ret <= pkg_stdLogicVector("01101001");
      when "11100101" =>
        zz_io_ret <= pkg_stdLogicVector("11011001");
      when "11100110" =>
        zz_io_ret <= pkg_stdLogicVector("10001110");
      when "11100111" =>
        zz_io_ret <= pkg_stdLogicVector("10010100");
      when "11101000" =>
        zz_io_ret <= pkg_stdLogicVector("10011011");
      when "11101001" =>
        zz_io_ret <= pkg_stdLogicVector("00011110");
      when "11101010" =>
        zz_io_ret <= pkg_stdLogicVector("10000111");
      when "11101011" =>
        zz_io_ret <= pkg_stdLogicVector("11101001");
      when "11101100" =>
        zz_io_ret <= pkg_stdLogicVector("11001110");
      when "11101101" =>
        zz_io_ret <= pkg_stdLogicVector("01010101");
      when "11101110" =>
        zz_io_ret <= pkg_stdLogicVector("00101000");
      when "11101111" =>
        zz_io_ret <= pkg_stdLogicVector("11011111");
      when "11110000" =>
        zz_io_ret <= pkg_stdLogicVector("10001100");
      when "11110001" =>
        zz_io_ret <= pkg_stdLogicVector("10100001");
      when "11110010" =>
        zz_io_ret <= pkg_stdLogicVector("10001001");
      when "11110011" =>
        zz_io_ret <= pkg_stdLogicVector("00001101");
      when "11110100" =>
        zz_io_ret <= pkg_stdLogicVector("10111111");
      when "11110101" =>
        zz_io_ret <= pkg_stdLogicVector("11100110");
      when "11110110" =>
        zz_io_ret <= pkg_stdLogicVector("01000010");
      when "11110111" =>
        zz_io_ret <= pkg_stdLogicVector("01101000");
      when "11111000" =>
        zz_io_ret <= pkg_stdLogicVector("01000001");
      when "11111001" =>
        zz_io_ret <= pkg_stdLogicVector("10011001");
      when "11111010" =>
        zz_io_ret <= pkg_stdLogicVector("00101101");
      when "11111011" =>
        zz_io_ret <= pkg_stdLogicVector("00001111");
      when "11111100" =>
        zz_io_ret <= pkg_stdLogicVector("10110000");
      when "11111101" =>
        zz_io_ret <= pkg_stdLogicVector("01010100");
      when "11111110" =>
        zz_io_ret <= pkg_stdLogicVector("10111011");
      when others =>
        zz_io_ret <= pkg_stdLogicVector("00010110");
    end case;
  end process;

  io_ret <= zz_io_ret;
end arch;


--SubByte_1 replaced by SubByte


--SubByte_2 replaced by SubByte


--SubByte_3 replaced by SubByte


--SubByte_4 replaced by SubByte


--SubByte_5 replaced by SubByte


--SubByte_6 replaced by SubByte


--SubByte_7 replaced by SubByte


--SubByte_8 replaced by SubByte


--SubByte_9 replaced by SubByte


--SubByte_10 replaced by SubByte


--SubByte_11 replaced by SubByte


--SubByte_12 replaced by SubByte


--SubByte_13 replaced by SubByte


--SubByte_14 replaced by SubByte


--SubByte_15 replaced by SubByte


--SubByte_16 replaced by SubByte


--SubByte_17 replaced by SubByte


--SubByte_18 replaced by SubByte


--SubByte_19 replaced by SubByte


--SubByte_20 replaced by SubByte


--SubByte_21 replaced by SubByte


--SubByte_22 replaced by SubByte


--SubByte_23 replaced by SubByte


--SubByte_24 replaced by SubByte


--SubByte_25 replaced by SubByte


--SubByte_26 replaced by SubByte


--SubByte_27 replaced by SubByte


--SubByte_28 replaced by SubByte


--SubByte_29 replaced by SubByte


--SubByte_30 replaced by SubByte


--SubByte_31 replaced by SubByte


--SubByte_32 replaced by SubByte


--SubByte_33 replaced by SubByte


--SubByte_34 replaced by SubByte


--SubByte_35 replaced by SubByte


--SubByte_36 replaced by SubByte


--SubByte_37 replaced by SubByte


--SubByte_38 replaced by SubByte


--SubByte_39 replaced by SubByte

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity SubWord is
  port(
    io_bs_0 : in std_logic_vector(7 downto 0);
    io_bs_1 : in std_logic_vector(7 downto 0);
    io_bs_2 : in std_logic_vector(7 downto 0);
    io_bs_3 : in std_logic_vector(7 downto 0);
    io_ret_0 : out std_logic_vector(7 downto 0);
    io_ret_1 : out std_logic_vector(7 downto 0);
    io_ret_2 : out std_logic_vector(7 downto 0);
    io_ret_3 : out std_logic_vector(7 downto 0)
  );
end SubWord;

architecture arch of SubWord is
  signal subByte_200_io_ret : std_logic_vector(7 downto 0);
  signal subByte_201_io_ret : std_logic_vector(7 downto 0);
  signal subByte_202_io_ret : std_logic_vector(7 downto 0);
  signal subByte_203_io_ret : std_logic_vector(7 downto 0);

begin
  subByte_200 : entity work.SubByte
    port map ( 
      io_b => io_bs_0,
      io_ret => subByte_200_io_ret 
    );
  subByte_201 : entity work.SubByte
    port map ( 
      io_b => io_bs_1,
      io_ret => subByte_201_io_ret 
    );
  subByte_202 : entity work.SubByte
    port map ( 
      io_b => io_bs_2,
      io_ret => subByte_202_io_ret 
    );
  subByte_203 : entity work.SubByte
    port map ( 
      io_b => io_bs_3,
      io_ret => subByte_203_io_ret 
    );
  io_ret_0 <= subByte_200_io_ret;
  io_ret_1 <= subByte_201_io_ret;
  io_ret_2 <= subByte_202_io_ret;
  io_ret_3 <= subByte_203_io_ret;
end arch;


--SubByte_40 replaced by SubByte


--SubByte_41 replaced by SubByte


--SubByte_42 replaced by SubByte


--SubByte_43 replaced by SubByte


--SubByte_44 replaced by SubByte


--SubByte_45 replaced by SubByte


--SubByte_46 replaced by SubByte


--SubByte_47 replaced by SubByte


--SubByte_48 replaced by SubByte


--SubByte_49 replaced by SubByte


--SubByte_50 replaced by SubByte


--SubByte_51 replaced by SubByte


--SubByte_52 replaced by SubByte


--SubByte_53 replaced by SubByte


--SubByte_54 replaced by SubByte


--SubByte_55 replaced by SubByte

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity MixColumn is
  port(
    io_c_0 : in std_logic_vector(7 downto 0);
    io_c_1 : in std_logic_vector(7 downto 0);
    io_c_2 : in std_logic_vector(7 downto 0);
    io_c_3 : in std_logic_vector(7 downto 0);
    io_ret_0 : out std_logic_vector(7 downto 0);
    io_ret_1 : out std_logic_vector(7 downto 0);
    io_ret_2 : out std_logic_vector(7 downto 0);
    io_ret_3 : out std_logic_vector(7 downto 0)
  );
end MixColumn;

architecture arch of MixColumn is

  signal zz_io_ret_0 : std_logic_vector(7 downto 0);
  signal when_AES_Round_l160 : std_logic;
  signal zz_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal when_AES_Round_l160_1 : std_logic;
  signal zz_io_ret_1 : std_logic_vector(7 downto 0);
  signal when_AES_Round_l160_2 : std_logic;
  signal zz_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal when_AES_Round_l160_3 : std_logic;
  signal zz_io_ret_2 : std_logic_vector(7 downto 0);
  signal when_AES_Round_l160_4 : std_logic;
  signal zz_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal when_AES_Round_l160_5 : std_logic;
  signal zz_io_ret_3 : std_logic_vector(7 downto 0);
  signal when_AES_Round_l160_6 : std_logic;
  signal zz_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal when_AES_Round_l160_7 : std_logic;
begin
  when_AES_Round_l160 <= pkg_toStdLogic(pkg_extract(io_c_0,7) = pkg_toStdLogic(false));
  process(when_AES_Round_l160,io_c_0)
  begin
    if when_AES_Round_l160 = '1' then
      zz_io_ret_0 <= std_logic_vector(shift_left(unsigned(io_c_0),1));
    else
      zz_io_ret_0 <= (std_logic_vector(shift_left(unsigned(io_c_0),1)) xor pkg_stdLogicVector("00011011"));
    end if;
  end process;

  when_AES_Round_l160_1 <= pkg_toStdLogic(pkg_extract(io_c_1,7) = pkg_toStdLogic(false));
  process(when_AES_Round_l160_1,io_c_1)
  begin
    if when_AES_Round_l160_1 = '1' then
      zz_io_ret_0_1 <= std_logic_vector(shift_left(unsigned(io_c_1),1));
    else
      zz_io_ret_0_1 <= (std_logic_vector(shift_left(unsigned(io_c_1),1)) xor pkg_stdLogicVector("00011011"));
    end if;
  end process;

  io_ret_0 <= (((zz_io_ret_0 xor (zz_io_ret_0_1 xor io_c_1)) xor io_c_2) xor io_c_3);
  when_AES_Round_l160_2 <= pkg_toStdLogic(pkg_extract(io_c_1,7) = pkg_toStdLogic(false));
  process(when_AES_Round_l160_2,io_c_1)
  begin
    if when_AES_Round_l160_2 = '1' then
      zz_io_ret_1 <= std_logic_vector(shift_left(unsigned(io_c_1),1));
    else
      zz_io_ret_1 <= (std_logic_vector(shift_left(unsigned(io_c_1),1)) xor pkg_stdLogicVector("00011011"));
    end if;
  end process;

  when_AES_Round_l160_3 <= pkg_toStdLogic(pkg_extract(io_c_2,7) = pkg_toStdLogic(false));
  process(when_AES_Round_l160_3,io_c_2)
  begin
    if when_AES_Round_l160_3 = '1' then
      zz_io_ret_1_1 <= std_logic_vector(shift_left(unsigned(io_c_2),1));
    else
      zz_io_ret_1_1 <= (std_logic_vector(shift_left(unsigned(io_c_2),1)) xor pkg_stdLogicVector("00011011"));
    end if;
  end process;

  io_ret_1 <= (((io_c_0 xor zz_io_ret_1) xor (zz_io_ret_1_1 xor io_c_2)) xor io_c_3);
  when_AES_Round_l160_4 <= pkg_toStdLogic(pkg_extract(io_c_2,7) = pkg_toStdLogic(false));
  process(when_AES_Round_l160_4,io_c_2)
  begin
    if when_AES_Round_l160_4 = '1' then
      zz_io_ret_2 <= std_logic_vector(shift_left(unsigned(io_c_2),1));
    else
      zz_io_ret_2 <= (std_logic_vector(shift_left(unsigned(io_c_2),1)) xor pkg_stdLogicVector("00011011"));
    end if;
  end process;

  when_AES_Round_l160_5 <= pkg_toStdLogic(pkg_extract(io_c_3,7) = pkg_toStdLogic(false));
  process(when_AES_Round_l160_5,io_c_3)
  begin
    if when_AES_Round_l160_5 = '1' then
      zz_io_ret_2_1 <= std_logic_vector(shift_left(unsigned(io_c_3),1));
    else
      zz_io_ret_2_1 <= (std_logic_vector(shift_left(unsigned(io_c_3),1)) xor pkg_stdLogicVector("00011011"));
    end if;
  end process;

  io_ret_2 <= (((io_c_0 xor io_c_1) xor zz_io_ret_2) xor (zz_io_ret_2_1 xor io_c_3));
  when_AES_Round_l160_6 <= pkg_toStdLogic(pkg_extract(io_c_0,7) = pkg_toStdLogic(false));
  process(when_AES_Round_l160_6,io_c_0)
  begin
    if when_AES_Round_l160_6 = '1' then
      zz_io_ret_3 <= std_logic_vector(shift_left(unsigned(io_c_0),1));
    else
      zz_io_ret_3 <= (std_logic_vector(shift_left(unsigned(io_c_0),1)) xor pkg_stdLogicVector("00011011"));
    end if;
  end process;

  when_AES_Round_l160_7 <= pkg_toStdLogic(pkg_extract(io_c_3,7) = pkg_toStdLogic(false));
  process(when_AES_Round_l160_7,io_c_3)
  begin
    if when_AES_Round_l160_7 = '1' then
      zz_io_ret_3_1 <= std_logic_vector(shift_left(unsigned(io_c_3),1));
    else
      zz_io_ret_3_1 <= (std_logic_vector(shift_left(unsigned(io_c_3),1)) xor pkg_stdLogicVector("00011011"));
    end if;
  end process;

  io_ret_3 <= ((((zz_io_ret_3 xor io_c_0) xor io_c_1) xor io_c_2) xor zz_io_ret_3_1);
end arch;


--MixColumn_1 replaced by MixColumn


--MixColumn_2 replaced by MixColumn


--MixColumn_3 replaced by MixColumn


--SubWord_1 replaced by SubWord


--SubByte_56 replaced by SubByte


--SubByte_57 replaced by SubByte


--SubByte_58 replaced by SubByte


--SubByte_59 replaced by SubByte


--SubByte_60 replaced by SubByte


--SubByte_61 replaced by SubByte


--SubByte_62 replaced by SubByte


--SubByte_63 replaced by SubByte


--SubByte_64 replaced by SubByte


--SubByte_65 replaced by SubByte


--SubByte_66 replaced by SubByte


--SubByte_67 replaced by SubByte


--SubByte_68 replaced by SubByte


--SubByte_69 replaced by SubByte


--SubByte_70 replaced by SubByte


--SubByte_71 replaced by SubByte


--MixColumn_4 replaced by MixColumn


--MixColumn_5 replaced by MixColumn


--MixColumn_6 replaced by MixColumn


--MixColumn_7 replaced by MixColumn


--SubWord_2 replaced by SubWord


--SubByte_72 replaced by SubByte


--SubByte_73 replaced by SubByte


--SubByte_74 replaced by SubByte


--SubByte_75 replaced by SubByte


--SubByte_76 replaced by SubByte


--SubByte_77 replaced by SubByte


--SubByte_78 replaced by SubByte


--SubByte_79 replaced by SubByte


--SubByte_80 replaced by SubByte


--SubByte_81 replaced by SubByte


--SubByte_82 replaced by SubByte


--SubByte_83 replaced by SubByte


--SubByte_84 replaced by SubByte


--SubByte_85 replaced by SubByte


--SubByte_86 replaced by SubByte


--SubByte_87 replaced by SubByte


--MixColumn_8 replaced by MixColumn


--MixColumn_9 replaced by MixColumn


--MixColumn_10 replaced by MixColumn


--MixColumn_11 replaced by MixColumn


--SubWord_3 replaced by SubWord


--SubByte_88 replaced by SubByte


--SubByte_89 replaced by SubByte


--SubByte_90 replaced by SubByte


--SubByte_91 replaced by SubByte


--SubByte_92 replaced by SubByte


--SubByte_93 replaced by SubByte


--SubByte_94 replaced by SubByte


--SubByte_95 replaced by SubByte


--SubByte_96 replaced by SubByte


--SubByte_97 replaced by SubByte


--SubByte_98 replaced by SubByte


--SubByte_99 replaced by SubByte


--SubByte_100 replaced by SubByte


--SubByte_101 replaced by SubByte


--SubByte_102 replaced by SubByte


--SubByte_103 replaced by SubByte


--MixColumn_12 replaced by MixColumn


--MixColumn_13 replaced by MixColumn


--MixColumn_14 replaced by MixColumn


--MixColumn_15 replaced by MixColumn


--SubWord_4 replaced by SubWord


--SubByte_104 replaced by SubByte


--SubByte_105 replaced by SubByte


--SubByte_106 replaced by SubByte


--SubByte_107 replaced by SubByte


--SubByte_108 replaced by SubByte


--SubByte_109 replaced by SubByte


--SubByte_110 replaced by SubByte


--SubByte_111 replaced by SubByte


--SubByte_112 replaced by SubByte


--SubByte_113 replaced by SubByte


--SubByte_114 replaced by SubByte


--SubByte_115 replaced by SubByte


--SubByte_116 replaced by SubByte


--SubByte_117 replaced by SubByte


--SubByte_118 replaced by SubByte


--SubByte_119 replaced by SubByte


--MixColumn_16 replaced by MixColumn


--MixColumn_17 replaced by MixColumn


--MixColumn_18 replaced by MixColumn


--MixColumn_19 replaced by MixColumn


--SubWord_5 replaced by SubWord


--SubByte_120 replaced by SubByte


--SubByte_121 replaced by SubByte


--SubByte_122 replaced by SubByte


--SubByte_123 replaced by SubByte


--SubByte_124 replaced by SubByte


--SubByte_125 replaced by SubByte


--SubByte_126 replaced by SubByte


--SubByte_127 replaced by SubByte


--SubByte_128 replaced by SubByte


--SubByte_129 replaced by SubByte


--SubByte_130 replaced by SubByte


--SubByte_131 replaced by SubByte


--SubByte_132 replaced by SubByte


--SubByte_133 replaced by SubByte


--SubByte_134 replaced by SubByte


--SubByte_135 replaced by SubByte


--MixColumn_20 replaced by MixColumn


--MixColumn_21 replaced by MixColumn


--MixColumn_22 replaced by MixColumn


--MixColumn_23 replaced by MixColumn


--SubWord_6 replaced by SubWord


--SubByte_136 replaced by SubByte


--SubByte_137 replaced by SubByte


--SubByte_138 replaced by SubByte


--SubByte_139 replaced by SubByte


--SubByte_140 replaced by SubByte


--SubByte_141 replaced by SubByte


--SubByte_142 replaced by SubByte


--SubByte_143 replaced by SubByte


--SubByte_144 replaced by SubByte


--SubByte_145 replaced by SubByte


--SubByte_146 replaced by SubByte


--SubByte_147 replaced by SubByte


--SubByte_148 replaced by SubByte


--SubByte_149 replaced by SubByte


--SubByte_150 replaced by SubByte


--SubByte_151 replaced by SubByte


--MixColumn_24 replaced by MixColumn


--MixColumn_25 replaced by MixColumn


--MixColumn_26 replaced by MixColumn


--MixColumn_27 replaced by MixColumn


--SubWord_7 replaced by SubWord


--SubByte_152 replaced by SubByte


--SubByte_153 replaced by SubByte


--SubByte_154 replaced by SubByte


--SubByte_155 replaced by SubByte


--SubByte_156 replaced by SubByte


--SubByte_157 replaced by SubByte


--SubByte_158 replaced by SubByte


--SubByte_159 replaced by SubByte


--SubByte_160 replaced by SubByte


--SubByte_161 replaced by SubByte


--SubByte_162 replaced by SubByte


--SubByte_163 replaced by SubByte


--SubByte_164 replaced by SubByte


--SubByte_165 replaced by SubByte


--SubByte_166 replaced by SubByte


--SubByte_167 replaced by SubByte


--MixColumn_28 replaced by MixColumn


--MixColumn_29 replaced by MixColumn


--MixColumn_30 replaced by MixColumn


--MixColumn_31 replaced by MixColumn


--SubWord_8 replaced by SubWord


--SubByte_168 replaced by SubByte


--SubByte_169 replaced by SubByte


--SubByte_170 replaced by SubByte


--SubByte_171 replaced by SubByte


--SubByte_172 replaced by SubByte


--SubByte_173 replaced by SubByte


--SubByte_174 replaced by SubByte


--SubByte_175 replaced by SubByte


--SubByte_176 replaced by SubByte


--SubByte_177 replaced by SubByte


--SubByte_178 replaced by SubByte


--SubByte_179 replaced by SubByte


--SubByte_180 replaced by SubByte


--SubByte_181 replaced by SubByte


--SubByte_182 replaced by SubByte


--SubByte_183 replaced by SubByte


--MixColumn_32 replaced by MixColumn


--MixColumn_33 replaced by MixColumn


--MixColumn_34 replaced by MixColumn


--MixColumn_35 replaced by MixColumn


--SubWord_9 replaced by SubWord


--SubByte_184 replaced by SubByte


--SubByte_185 replaced by SubByte


--SubByte_186 replaced by SubByte


--SubByte_187 replaced by SubByte


--SubByte_188 replaced by SubByte


--SubByte_189 replaced by SubByte


--SubByte_190 replaced by SubByte


--SubByte_191 replaced by SubByte


--SubByte_192 replaced by SubByte


--SubByte_193 replaced by SubByte


--SubByte_194 replaced by SubByte


--SubByte_195 replaced by SubByte


--SubByte_196 replaced by SubByte


--SubByte_197 replaced by SubByte


--SubByte_198 replaced by SubByte


--SubByte_199 replaced by SubByte

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity AddRoundKey is
  port(
    io_rk_0_0 : in std_logic_vector(7 downto 0);
    io_rk_0_1 : in std_logic_vector(7 downto 0);
    io_rk_0_2 : in std_logic_vector(7 downto 0);
    io_rk_0_3 : in std_logic_vector(7 downto 0);
    io_rk_1_0 : in std_logic_vector(7 downto 0);
    io_rk_1_1 : in std_logic_vector(7 downto 0);
    io_rk_1_2 : in std_logic_vector(7 downto 0);
    io_rk_1_3 : in std_logic_vector(7 downto 0);
    io_rk_2_0 : in std_logic_vector(7 downto 0);
    io_rk_2_1 : in std_logic_vector(7 downto 0);
    io_rk_2_2 : in std_logic_vector(7 downto 0);
    io_rk_2_3 : in std_logic_vector(7 downto 0);
    io_rk_3_0 : in std_logic_vector(7 downto 0);
    io_rk_3_1 : in std_logic_vector(7 downto 0);
    io_rk_3_2 : in std_logic_vector(7 downto 0);
    io_rk_3_3 : in std_logic_vector(7 downto 0);
    io_s_0_0 : in std_logic_vector(7 downto 0);
    io_s_0_1 : in std_logic_vector(7 downto 0);
    io_s_0_2 : in std_logic_vector(7 downto 0);
    io_s_0_3 : in std_logic_vector(7 downto 0);
    io_s_1_0 : in std_logic_vector(7 downto 0);
    io_s_1_1 : in std_logic_vector(7 downto 0);
    io_s_1_2 : in std_logic_vector(7 downto 0);
    io_s_1_3 : in std_logic_vector(7 downto 0);
    io_s_2_0 : in std_logic_vector(7 downto 0);
    io_s_2_1 : in std_logic_vector(7 downto 0);
    io_s_2_2 : in std_logic_vector(7 downto 0);
    io_s_2_3 : in std_logic_vector(7 downto 0);
    io_s_3_0 : in std_logic_vector(7 downto 0);
    io_s_3_1 : in std_logic_vector(7 downto 0);
    io_s_3_2 : in std_logic_vector(7 downto 0);
    io_s_3_3 : in std_logic_vector(7 downto 0);
    io_ret_0_0 : out std_logic_vector(7 downto 0);
    io_ret_0_1 : out std_logic_vector(7 downto 0);
    io_ret_0_2 : out std_logic_vector(7 downto 0);
    io_ret_0_3 : out std_logic_vector(7 downto 0);
    io_ret_1_0 : out std_logic_vector(7 downto 0);
    io_ret_1_1 : out std_logic_vector(7 downto 0);
    io_ret_1_2 : out std_logic_vector(7 downto 0);
    io_ret_1_3 : out std_logic_vector(7 downto 0);
    io_ret_2_0 : out std_logic_vector(7 downto 0);
    io_ret_2_1 : out std_logic_vector(7 downto 0);
    io_ret_2_2 : out std_logic_vector(7 downto 0);
    io_ret_2_3 : out std_logic_vector(7 downto 0);
    io_ret_3_0 : out std_logic_vector(7 downto 0);
    io_ret_3_1 : out std_logic_vector(7 downto 0);
    io_ret_3_2 : out std_logic_vector(7 downto 0);
    io_ret_3_3 : out std_logic_vector(7 downto 0)
  );
end AddRoundKey;

architecture arch of AddRoundKey is

begin
  io_ret_0_0 <= (io_rk_0_0 xor io_s_0_0);
  io_ret_0_1 <= (io_rk_0_1 xor io_s_0_1);
  io_ret_0_2 <= (io_rk_0_2 xor io_s_0_2);
  io_ret_0_3 <= (io_rk_0_3 xor io_s_0_3);
  io_ret_1_0 <= (io_rk_1_0 xor io_s_1_0);
  io_ret_1_1 <= (io_rk_1_1 xor io_s_1_1);
  io_ret_1_2 <= (io_rk_1_2 xor io_s_1_2);
  io_ret_1_3 <= (io_rk_1_3 xor io_s_1_3);
  io_ret_2_0 <= (io_rk_2_0 xor io_s_2_0);
  io_ret_2_1 <= (io_rk_2_1 xor io_s_2_1);
  io_ret_2_2 <= (io_rk_2_2 xor io_s_2_2);
  io_ret_2_3 <= (io_rk_2_3 xor io_s_2_3);
  io_ret_3_0 <= (io_rk_3_0 xor io_s_3_0);
  io_ret_3_1 <= (io_rk_3_1 xor io_s_3_1);
  io_ret_3_2 <= (io_rk_3_2 xor io_s_3_2);
  io_ret_3_3 <= (io_rk_3_3 xor io_s_3_3);
end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity NextRC is
  port(
    io_rc : in std_logic_vector(7 downto 0);
    io_ret : out std_logic_vector(7 downto 0)
  );
end NextRC;

architecture arch of NextRC is

  signal when_AES_Round_l199 : std_logic;
begin
  when_AES_Round_l199 <= pkg_toStdLogic(pkg_extract(io_rc,7) = pkg_toStdLogic(false));
  process(when_AES_Round_l199,io_rc)
  begin
    if when_AES_Round_l199 = '1' then
      io_ret <= std_logic_vector(shift_left(unsigned(io_rc),1));
    else
      io_ret <= (std_logic_vector(shift_left(unsigned(io_rc),1)) xor pkg_stdLogicVector("00011011"));
    end if;
  end process;

end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity KeySchedule is
  port(
    io_key_0_0 : in std_logic_vector(7 downto 0);
    io_key_0_1 : in std_logic_vector(7 downto 0);
    io_key_0_2 : in std_logic_vector(7 downto 0);
    io_key_0_3 : in std_logic_vector(7 downto 0);
    io_key_1_0 : in std_logic_vector(7 downto 0);
    io_key_1_1 : in std_logic_vector(7 downto 0);
    io_key_1_2 : in std_logic_vector(7 downto 0);
    io_key_1_3 : in std_logic_vector(7 downto 0);
    io_key_2_0 : in std_logic_vector(7 downto 0);
    io_key_2_1 : in std_logic_vector(7 downto 0);
    io_key_2_2 : in std_logic_vector(7 downto 0);
    io_key_2_3 : in std_logic_vector(7 downto 0);
    io_key_3_0 : in std_logic_vector(7 downto 0);
    io_key_3_1 : in std_logic_vector(7 downto 0);
    io_key_3_2 : in std_logic_vector(7 downto 0);
    io_key_3_3 : in std_logic_vector(7 downto 0);
    io_c : in std_logic_vector(7 downto 0);
    io_ret_0_0 : out std_logic_vector(7 downto 0);
    io_ret_0_1 : out std_logic_vector(7 downto 0);
    io_ret_0_2 : out std_logic_vector(7 downto 0);
    io_ret_0_3 : out std_logic_vector(7 downto 0);
    io_ret_1_0 : out std_logic_vector(7 downto 0);
    io_ret_1_1 : out std_logic_vector(7 downto 0);
    io_ret_1_2 : out std_logic_vector(7 downto 0);
    io_ret_1_3 : out std_logic_vector(7 downto 0);
    io_ret_2_0 : out std_logic_vector(7 downto 0);
    io_ret_2_1 : out std_logic_vector(7 downto 0);
    io_ret_2_2 : out std_logic_vector(7 downto 0);
    io_ret_2_3 : out std_logic_vector(7 downto 0);
    io_ret_3_0 : out std_logic_vector(7 downto 0);
    io_ret_3_1 : out std_logic_vector(7 downto 0);
    io_ret_3_2 : out std_logic_vector(7 downto 0);
    io_ret_3_3 : out std_logic_vector(7 downto 0)
  );
end KeySchedule;

architecture arch of KeySchedule is
  signal subword_10_io_ret_0 : std_logic_vector(7 downto 0);
  signal subword_10_io_ret_1 : std_logic_vector(7 downto 0);
  signal subword_10_io_ret_2 : std_logic_vector(7 downto 0);
  signal subword_10_io_ret_3 : std_logic_vector(7 downto 0);

  signal keyT_0_0 : std_logic_vector(7 downto 0);
  signal keyT_0_1 : std_logic_vector(7 downto 0);
  signal keyT_0_2 : std_logic_vector(7 downto 0);
  signal keyT_0_3 : std_logic_vector(7 downto 0);
  signal keyT_1_0 : std_logic_vector(7 downto 0);
  signal keyT_1_1 : std_logic_vector(7 downto 0);
  signal keyT_1_2 : std_logic_vector(7 downto 0);
  signal keyT_1_3 : std_logic_vector(7 downto 0);
  signal keyT_2_0 : std_logic_vector(7 downto 0);
  signal keyT_2_1 : std_logic_vector(7 downto 0);
  signal keyT_2_2 : std_logic_vector(7 downto 0);
  signal keyT_2_3 : std_logic_vector(7 downto 0);
  signal keyT_3_0 : std_logic_vector(7 downto 0);
  signal keyT_3_1 : std_logic_vector(7 downto 0);
  signal keyT_3_2 : std_logic_vector(7 downto 0);
  signal keyT_3_3 : std_logic_vector(7 downto 0);
  signal w0_0 : std_logic_vector(7 downto 0);
  signal w0_1 : std_logic_vector(7 downto 0);
  signal w0_2 : std_logic_vector(7 downto 0);
  signal w0_3 : std_logic_vector(7 downto 0);
  signal w1_0 : std_logic_vector(7 downto 0);
  signal w1_1 : std_logic_vector(7 downto 0);
  signal w1_2 : std_logic_vector(7 downto 0);
  signal w1_3 : std_logic_vector(7 downto 0);
  signal w2_0 : std_logic_vector(7 downto 0);
  signal w2_1 : std_logic_vector(7 downto 0);
  signal w2_2 : std_logic_vector(7 downto 0);
  signal w2_3 : std_logic_vector(7 downto 0);
  signal w3_0 : std_logic_vector(7 downto 0);
  signal w3_1 : std_logic_vector(7 downto 0);
  signal w3_2 : std_logic_vector(7 downto 0);
  signal w3_3 : std_logic_vector(7 downto 0);
begin
  subword_10 : entity work.SubWord
    port map ( 
      io_bs_0 => keyT_3_0,
      io_bs_1 => keyT_3_1,
      io_bs_2 => keyT_3_2,
      io_bs_3 => keyT_3_3,
      io_ret_0 => subword_10_io_ret_0,
      io_ret_1 => subword_10_io_ret_1,
      io_ret_2 => subword_10_io_ret_2,
      io_ret_3 => subword_10_io_ret_3 
    );
  keyT_0_0 <= io_key_0_0;
  keyT_0_1 <= io_key_1_0;
  keyT_0_2 <= io_key_2_0;
  keyT_0_3 <= io_key_3_0;
  keyT_1_0 <= io_key_0_1;
  keyT_1_1 <= io_key_1_1;
  keyT_1_2 <= io_key_2_1;
  keyT_1_3 <= io_key_3_1;
  keyT_2_0 <= io_key_0_2;
  keyT_2_1 <= io_key_1_2;
  keyT_2_2 <= io_key_2_2;
  keyT_2_3 <= io_key_3_2;
  keyT_3_0 <= io_key_0_3;
  keyT_3_1 <= io_key_1_3;
  keyT_3_2 <= io_key_2_3;
  keyT_3_3 <= io_key_3_3;
  w0_0 <= ((keyT_0_0 xor subword_10_io_ret_1) xor io_c);
  w0_1 <= ((keyT_0_1 xor subword_10_io_ret_2) xor pkg_stdLogicVector("00000000"));
  w0_2 <= ((keyT_0_2 xor subword_10_io_ret_3) xor pkg_stdLogicVector("00000000"));
  w0_3 <= ((keyT_0_3 xor subword_10_io_ret_0) xor pkg_stdLogicVector("00000000"));
  w1_0 <= (keyT_1_0 xor w0_0);
  w1_1 <= (keyT_1_1 xor w0_1);
  w1_2 <= (keyT_1_2 xor w0_2);
  w1_3 <= (keyT_1_3 xor w0_3);
  w2_0 <= (keyT_2_0 xor w1_0);
  w2_1 <= (keyT_2_1 xor w1_1);
  w2_2 <= (keyT_2_2 xor w1_2);
  w2_3 <= (keyT_2_3 xor w1_3);
  w3_0 <= (keyT_3_0 xor w2_0);
  w3_1 <= (keyT_3_1 xor w2_1);
  w3_2 <= (keyT_3_2 xor w2_2);
  w3_3 <= (keyT_3_3 xor w2_3);
  io_ret_0_0 <= w0_0;
  io_ret_0_1 <= w1_0;
  io_ret_0_2 <= w2_0;
  io_ret_0_3 <= w3_0;
  io_ret_1_0 <= w0_1;
  io_ret_1_1 <= w1_1;
  io_ret_1_2 <= w2_1;
  io_ret_1_3 <= w3_1;
  io_ret_2_0 <= w0_2;
  io_ret_2_1 <= w1_2;
  io_ret_2_2 <= w2_2;
  io_ret_2_3 <= w3_2;
  io_ret_3_0 <= w0_3;
  io_ret_3_1 <= w1_3;
  io_ret_3_2 <= w2_3;
  io_ret_3_3 <= w3_3;
end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity SubBytes is
  port(
    io_state_0_0 : in std_logic_vector(7 downto 0);
    io_state_0_1 : in std_logic_vector(7 downto 0);
    io_state_0_2 : in std_logic_vector(7 downto 0);
    io_state_0_3 : in std_logic_vector(7 downto 0);
    io_state_1_0 : in std_logic_vector(7 downto 0);
    io_state_1_1 : in std_logic_vector(7 downto 0);
    io_state_1_2 : in std_logic_vector(7 downto 0);
    io_state_1_3 : in std_logic_vector(7 downto 0);
    io_state_2_0 : in std_logic_vector(7 downto 0);
    io_state_2_1 : in std_logic_vector(7 downto 0);
    io_state_2_2 : in std_logic_vector(7 downto 0);
    io_state_2_3 : in std_logic_vector(7 downto 0);
    io_state_3_0 : in std_logic_vector(7 downto 0);
    io_state_3_1 : in std_logic_vector(7 downto 0);
    io_state_3_2 : in std_logic_vector(7 downto 0);
    io_state_3_3 : in std_logic_vector(7 downto 0);
    io_ret_0_0 : out std_logic_vector(7 downto 0);
    io_ret_0_1 : out std_logic_vector(7 downto 0);
    io_ret_0_2 : out std_logic_vector(7 downto 0);
    io_ret_0_3 : out std_logic_vector(7 downto 0);
    io_ret_1_0 : out std_logic_vector(7 downto 0);
    io_ret_1_1 : out std_logic_vector(7 downto 0);
    io_ret_1_2 : out std_logic_vector(7 downto 0);
    io_ret_1_3 : out std_logic_vector(7 downto 0);
    io_ret_2_0 : out std_logic_vector(7 downto 0);
    io_ret_2_1 : out std_logic_vector(7 downto 0);
    io_ret_2_2 : out std_logic_vector(7 downto 0);
    io_ret_2_3 : out std_logic_vector(7 downto 0);
    io_ret_3_0 : out std_logic_vector(7 downto 0);
    io_ret_3_1 : out std_logic_vector(7 downto 0);
    io_ret_3_2 : out std_logic_vector(7 downto 0);
    io_ret_3_3 : out std_logic_vector(7 downto 0)
  );
end SubBytes;

architecture arch of SubBytes is
  signal subByte_200_io_ret : std_logic_vector(7 downto 0);
  signal subByte_201_io_ret : std_logic_vector(7 downto 0);
  signal subByte_202_io_ret : std_logic_vector(7 downto 0);
  signal subByte_203_io_ret : std_logic_vector(7 downto 0);
  signal subByte_204_io_ret : std_logic_vector(7 downto 0);
  signal subByte_205_io_ret : std_logic_vector(7 downto 0);
  signal subByte_206_io_ret : std_logic_vector(7 downto 0);
  signal subByte_207_io_ret : std_logic_vector(7 downto 0);
  signal subByte_208_io_ret : std_logic_vector(7 downto 0);
  signal subByte_209_io_ret : std_logic_vector(7 downto 0);
  signal subByte_210_io_ret : std_logic_vector(7 downto 0);
  signal subByte_211_io_ret : std_logic_vector(7 downto 0);
  signal subByte_212_io_ret : std_logic_vector(7 downto 0);
  signal subByte_213_io_ret : std_logic_vector(7 downto 0);
  signal subByte_214_io_ret : std_logic_vector(7 downto 0);
  signal subByte_215_io_ret : std_logic_vector(7 downto 0);

begin
  subByte_200 : entity work.SubByte
    port map ( 
      io_b => io_state_0_0,
      io_ret => subByte_200_io_ret 
    );
  subByte_201 : entity work.SubByte
    port map ( 
      io_b => io_state_0_1,
      io_ret => subByte_201_io_ret 
    );
  subByte_202 : entity work.SubByte
    port map ( 
      io_b => io_state_0_2,
      io_ret => subByte_202_io_ret 
    );
  subByte_203 : entity work.SubByte
    port map ( 
      io_b => io_state_0_3,
      io_ret => subByte_203_io_ret 
    );
  subByte_204 : entity work.SubByte
    port map ( 
      io_b => io_state_1_0,
      io_ret => subByte_204_io_ret 
    );
  subByte_205 : entity work.SubByte
    port map ( 
      io_b => io_state_1_1,
      io_ret => subByte_205_io_ret 
    );
  subByte_206 : entity work.SubByte
    port map ( 
      io_b => io_state_1_2,
      io_ret => subByte_206_io_ret 
    );
  subByte_207 : entity work.SubByte
    port map ( 
      io_b => io_state_1_3,
      io_ret => subByte_207_io_ret 
    );
  subByte_208 : entity work.SubByte
    port map ( 
      io_b => io_state_2_0,
      io_ret => subByte_208_io_ret 
    );
  subByte_209 : entity work.SubByte
    port map ( 
      io_b => io_state_2_1,
      io_ret => subByte_209_io_ret 
    );
  subByte_210 : entity work.SubByte
    port map ( 
      io_b => io_state_2_2,
      io_ret => subByte_210_io_ret 
    );
  subByte_211 : entity work.SubByte
    port map ( 
      io_b => io_state_2_3,
      io_ret => subByte_211_io_ret 
    );
  subByte_212 : entity work.SubByte
    port map ( 
      io_b => io_state_3_0,
      io_ret => subByte_212_io_ret 
    );
  subByte_213 : entity work.SubByte
    port map ( 
      io_b => io_state_3_1,
      io_ret => subByte_213_io_ret 
    );
  subByte_214 : entity work.SubByte
    port map ( 
      io_b => io_state_3_2,
      io_ret => subByte_214_io_ret 
    );
  subByte_215 : entity work.SubByte
    port map ( 
      io_b => io_state_3_3,
      io_ret => subByte_215_io_ret 
    );
  io_ret_0_0 <= subByte_200_io_ret;
  io_ret_0_1 <= subByte_201_io_ret;
  io_ret_0_2 <= subByte_202_io_ret;
  io_ret_0_3 <= subByte_203_io_ret;
  io_ret_1_0 <= subByte_204_io_ret;
  io_ret_1_1 <= subByte_205_io_ret;
  io_ret_1_2 <= subByte_206_io_ret;
  io_ret_1_3 <= subByte_207_io_ret;
  io_ret_2_0 <= subByte_208_io_ret;
  io_ret_2_1 <= subByte_209_io_ret;
  io_ret_2_2 <= subByte_210_io_ret;
  io_ret_2_3 <= subByte_211_io_ret;
  io_ret_3_0 <= subByte_212_io_ret;
  io_ret_3_1 <= subByte_213_io_ret;
  io_ret_3_2 <= subByte_214_io_ret;
  io_ret_3_3 <= subByte_215_io_ret;
end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity ShiftRows is
  port(
    io_state_0_0 : in std_logic_vector(7 downto 0);
    io_state_0_1 : in std_logic_vector(7 downto 0);
    io_state_0_2 : in std_logic_vector(7 downto 0);
    io_state_0_3 : in std_logic_vector(7 downto 0);
    io_state_1_0 : in std_logic_vector(7 downto 0);
    io_state_1_1 : in std_logic_vector(7 downto 0);
    io_state_1_2 : in std_logic_vector(7 downto 0);
    io_state_1_3 : in std_logic_vector(7 downto 0);
    io_state_2_0 : in std_logic_vector(7 downto 0);
    io_state_2_1 : in std_logic_vector(7 downto 0);
    io_state_2_2 : in std_logic_vector(7 downto 0);
    io_state_2_3 : in std_logic_vector(7 downto 0);
    io_state_3_0 : in std_logic_vector(7 downto 0);
    io_state_3_1 : in std_logic_vector(7 downto 0);
    io_state_3_2 : in std_logic_vector(7 downto 0);
    io_state_3_3 : in std_logic_vector(7 downto 0);
    io_ret_0_0 : out std_logic_vector(7 downto 0);
    io_ret_0_1 : out std_logic_vector(7 downto 0);
    io_ret_0_2 : out std_logic_vector(7 downto 0);
    io_ret_0_3 : out std_logic_vector(7 downto 0);
    io_ret_1_0 : out std_logic_vector(7 downto 0);
    io_ret_1_1 : out std_logic_vector(7 downto 0);
    io_ret_1_2 : out std_logic_vector(7 downto 0);
    io_ret_1_3 : out std_logic_vector(7 downto 0);
    io_ret_2_0 : out std_logic_vector(7 downto 0);
    io_ret_2_1 : out std_logic_vector(7 downto 0);
    io_ret_2_2 : out std_logic_vector(7 downto 0);
    io_ret_2_3 : out std_logic_vector(7 downto 0);
    io_ret_3_0 : out std_logic_vector(7 downto 0);
    io_ret_3_1 : out std_logic_vector(7 downto 0);
    io_ret_3_2 : out std_logic_vector(7 downto 0);
    io_ret_3_3 : out std_logic_vector(7 downto 0)
  );
end ShiftRows;

architecture arch of ShiftRows is

begin
  io_ret_0_0 <= io_state_0_0;
  io_ret_0_1 <= io_state_0_1;
  io_ret_0_2 <= io_state_0_2;
  io_ret_0_3 <= io_state_0_3;
  io_ret_1_0 <= io_state_1_1;
  io_ret_1_1 <= io_state_1_2;
  io_ret_1_2 <= io_state_1_3;
  io_ret_1_3 <= io_state_1_0;
  io_ret_2_0 <= io_state_2_2;
  io_ret_2_1 <= io_state_2_3;
  io_ret_2_2 <= io_state_2_0;
  io_ret_2_3 <= io_state_2_1;
  io_ret_3_0 <= io_state_3_3;
  io_ret_3_1 <= io_state_3_0;
  io_ret_3_2 <= io_state_3_1;
  io_ret_3_3 <= io_state_3_2;
end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity MixColumns is
  port(
    io_state_0_0 : in std_logic_vector(7 downto 0);
    io_state_0_1 : in std_logic_vector(7 downto 0);
    io_state_0_2 : in std_logic_vector(7 downto 0);
    io_state_0_3 : in std_logic_vector(7 downto 0);
    io_state_1_0 : in std_logic_vector(7 downto 0);
    io_state_1_1 : in std_logic_vector(7 downto 0);
    io_state_1_2 : in std_logic_vector(7 downto 0);
    io_state_1_3 : in std_logic_vector(7 downto 0);
    io_state_2_0 : in std_logic_vector(7 downto 0);
    io_state_2_1 : in std_logic_vector(7 downto 0);
    io_state_2_2 : in std_logic_vector(7 downto 0);
    io_state_2_3 : in std_logic_vector(7 downto 0);
    io_state_3_0 : in std_logic_vector(7 downto 0);
    io_state_3_1 : in std_logic_vector(7 downto 0);
    io_state_3_2 : in std_logic_vector(7 downto 0);
    io_state_3_3 : in std_logic_vector(7 downto 0);
    io_ret_0_0 : out std_logic_vector(7 downto 0);
    io_ret_0_1 : out std_logic_vector(7 downto 0);
    io_ret_0_2 : out std_logic_vector(7 downto 0);
    io_ret_0_3 : out std_logic_vector(7 downto 0);
    io_ret_1_0 : out std_logic_vector(7 downto 0);
    io_ret_1_1 : out std_logic_vector(7 downto 0);
    io_ret_1_2 : out std_logic_vector(7 downto 0);
    io_ret_1_3 : out std_logic_vector(7 downto 0);
    io_ret_2_0 : out std_logic_vector(7 downto 0);
    io_ret_2_1 : out std_logic_vector(7 downto 0);
    io_ret_2_2 : out std_logic_vector(7 downto 0);
    io_ret_2_3 : out std_logic_vector(7 downto 0);
    io_ret_3_0 : out std_logic_vector(7 downto 0);
    io_ret_3_1 : out std_logic_vector(7 downto 0);
    io_ret_3_2 : out std_logic_vector(7 downto 0);
    io_ret_3_3 : out std_logic_vector(7 downto 0)
  );
end MixColumns;

architecture arch of MixColumns is
  signal mixColumn_36_io_ret_0 : std_logic_vector(7 downto 0);
  signal mixColumn_36_io_ret_1 : std_logic_vector(7 downto 0);
  signal mixColumn_36_io_ret_2 : std_logic_vector(7 downto 0);
  signal mixColumn_36_io_ret_3 : std_logic_vector(7 downto 0);
  signal mixColumn_37_io_ret_0 : std_logic_vector(7 downto 0);
  signal mixColumn_37_io_ret_1 : std_logic_vector(7 downto 0);
  signal mixColumn_37_io_ret_2 : std_logic_vector(7 downto 0);
  signal mixColumn_37_io_ret_3 : std_logic_vector(7 downto 0);
  signal mixColumn_38_io_ret_0 : std_logic_vector(7 downto 0);
  signal mixColumn_38_io_ret_1 : std_logic_vector(7 downto 0);
  signal mixColumn_38_io_ret_2 : std_logic_vector(7 downto 0);
  signal mixColumn_38_io_ret_3 : std_logic_vector(7 downto 0);
  signal mixColumn_39_io_ret_0 : std_logic_vector(7 downto 0);
  signal mixColumn_39_io_ret_1 : std_logic_vector(7 downto 0);
  signal mixColumn_39_io_ret_2 : std_logic_vector(7 downto 0);
  signal mixColumn_39_io_ret_3 : std_logic_vector(7 downto 0);

  signal ret_0_0 : std_logic_vector(7 downto 0);
  signal ret_0_1 : std_logic_vector(7 downto 0);
  signal ret_0_2 : std_logic_vector(7 downto 0);
  signal ret_0_3 : std_logic_vector(7 downto 0);
  signal ret_1_0 : std_logic_vector(7 downto 0);
  signal ret_1_1 : std_logic_vector(7 downto 0);
  signal ret_1_2 : std_logic_vector(7 downto 0);
  signal ret_1_3 : std_logic_vector(7 downto 0);
  signal ret_2_0 : std_logic_vector(7 downto 0);
  signal ret_2_1 : std_logic_vector(7 downto 0);
  signal ret_2_2 : std_logic_vector(7 downto 0);
  signal ret_2_3 : std_logic_vector(7 downto 0);
  signal ret_3_0 : std_logic_vector(7 downto 0);
  signal ret_3_1 : std_logic_vector(7 downto 0);
  signal ret_3_2 : std_logic_vector(7 downto 0);
  signal ret_3_3 : std_logic_vector(7 downto 0);
begin
  mixColumn_36 : entity work.MixColumn
    port map ( 
      io_c_0 => io_state_0_0,
      io_c_1 => io_state_1_0,
      io_c_2 => io_state_2_0,
      io_c_3 => io_state_3_0,
      io_ret_0 => mixColumn_36_io_ret_0,
      io_ret_1 => mixColumn_36_io_ret_1,
      io_ret_2 => mixColumn_36_io_ret_2,
      io_ret_3 => mixColumn_36_io_ret_3 
    );
  mixColumn_37 : entity work.MixColumn
    port map ( 
      io_c_0 => io_state_0_1,
      io_c_1 => io_state_1_1,
      io_c_2 => io_state_2_1,
      io_c_3 => io_state_3_1,
      io_ret_0 => mixColumn_37_io_ret_0,
      io_ret_1 => mixColumn_37_io_ret_1,
      io_ret_2 => mixColumn_37_io_ret_2,
      io_ret_3 => mixColumn_37_io_ret_3 
    );
  mixColumn_38 : entity work.MixColumn
    port map ( 
      io_c_0 => io_state_0_2,
      io_c_1 => io_state_1_2,
      io_c_2 => io_state_2_2,
      io_c_3 => io_state_3_2,
      io_ret_0 => mixColumn_38_io_ret_0,
      io_ret_1 => mixColumn_38_io_ret_1,
      io_ret_2 => mixColumn_38_io_ret_2,
      io_ret_3 => mixColumn_38_io_ret_3 
    );
  mixColumn_39 : entity work.MixColumn
    port map ( 
      io_c_0 => io_state_0_3,
      io_c_1 => io_state_1_3,
      io_c_2 => io_state_2_3,
      io_c_3 => io_state_3_3,
      io_ret_0 => mixColumn_39_io_ret_0,
      io_ret_1 => mixColumn_39_io_ret_1,
      io_ret_2 => mixColumn_39_io_ret_2,
      io_ret_3 => mixColumn_39_io_ret_3 
    );
  ret_0_0 <= mixColumn_36_io_ret_0;
  ret_0_1 <= mixColumn_36_io_ret_1;
  ret_0_2 <= mixColumn_36_io_ret_2;
  ret_0_3 <= mixColumn_36_io_ret_3;
  ret_1_0 <= mixColumn_37_io_ret_0;
  ret_1_1 <= mixColumn_37_io_ret_1;
  ret_1_2 <= mixColumn_37_io_ret_2;
  ret_1_3 <= mixColumn_37_io_ret_3;
  ret_2_0 <= mixColumn_38_io_ret_0;
  ret_2_1 <= mixColumn_38_io_ret_1;
  ret_2_2 <= mixColumn_38_io_ret_2;
  ret_2_3 <= mixColumn_38_io_ret_3;
  ret_3_0 <= mixColumn_39_io_ret_0;
  ret_3_1 <= mixColumn_39_io_ret_1;
  ret_3_2 <= mixColumn_39_io_ret_2;
  ret_3_3 <= mixColumn_39_io_ret_3;
  io_ret_0_0 <= ret_0_0;
  io_ret_0_1 <= ret_1_0;
  io_ret_0_2 <= ret_2_0;
  io_ret_0_3 <= ret_3_0;
  io_ret_1_0 <= ret_0_1;
  io_ret_1_1 <= ret_1_1;
  io_ret_1_2 <= ret_2_1;
  io_ret_1_3 <= ret_3_1;
  io_ret_2_0 <= ret_0_2;
  io_ret_2_1 <= ret_1_2;
  io_ret_2_2 <= ret_2_2;
  io_ret_2_3 <= ret_3_2;
  io_ret_3_0 <= ret_0_3;
  io_ret_3_1 <= ret_1_3;
  io_ret_3_2 <= ret_2_3;
  io_ret_3_3 <= ret_3_3;
end arch;


--AddRoundKey_1 replaced by AddRoundKey


--NextRC_1 replaced by NextRC


--KeySchedule_1 replaced by KeySchedule


--SubBytes_1 replaced by SubBytes


--ShiftRows_1 replaced by ShiftRows


--MixColumns_1 replaced by MixColumns


--AddRoundKey_2 replaced by AddRoundKey


--NextRC_2 replaced by NextRC


--KeySchedule_2 replaced by KeySchedule


--SubBytes_2 replaced by SubBytes


--ShiftRows_2 replaced by ShiftRows


--MixColumns_2 replaced by MixColumns


--AddRoundKey_3 replaced by AddRoundKey


--NextRC_3 replaced by NextRC


--KeySchedule_3 replaced by KeySchedule


--SubBytes_3 replaced by SubBytes


--ShiftRows_3 replaced by ShiftRows


--MixColumns_3 replaced by MixColumns


--AddRoundKey_4 replaced by AddRoundKey


--NextRC_4 replaced by NextRC


--KeySchedule_4 replaced by KeySchedule


--SubBytes_4 replaced by SubBytes


--ShiftRows_4 replaced by ShiftRows


--MixColumns_4 replaced by MixColumns


--AddRoundKey_5 replaced by AddRoundKey


--NextRC_5 replaced by NextRC


--KeySchedule_5 replaced by KeySchedule


--SubBytes_5 replaced by SubBytes


--ShiftRows_5 replaced by ShiftRows


--MixColumns_5 replaced by MixColumns


--AddRoundKey_6 replaced by AddRoundKey


--NextRC_6 replaced by NextRC


--KeySchedule_6 replaced by KeySchedule


--SubBytes_6 replaced by SubBytes


--ShiftRows_6 replaced by ShiftRows


--MixColumns_6 replaced by MixColumns


--AddRoundKey_7 replaced by AddRoundKey


--NextRC_7 replaced by NextRC


--KeySchedule_7 replaced by KeySchedule


--SubBytes_7 replaced by SubBytes


--ShiftRows_7 replaced by ShiftRows


--MixColumns_7 replaced by MixColumns


--AddRoundKey_8 replaced by AddRoundKey


--NextRC_8 replaced by NextRC


--KeySchedule_8 replaced by KeySchedule


--SubBytes_8 replaced by SubBytes


--ShiftRows_8 replaced by ShiftRows


--MixColumns_8 replaced by MixColumns


--AddRoundKey_9 replaced by AddRoundKey


--NextRC_9 replaced by NextRC


--KeySchedule_9 replaced by KeySchedule


--SubBytes_9 replaced by SubBytes


--ShiftRows_9 replaced by ShiftRows


--AddRoundKey_10 replaced by AddRoundKey

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity aesEncrypt_Unrolled is
  port(
    io_pt : in std_logic_vector(127 downto 0);
    io_key : in std_logic_vector(127 downto 0);
    io_ret : out std_logic_vector(127 downto 0);
    clk : in std_logic;
    reset : in std_logic
  );
end aesEncrypt_Unrolled;

architecture arch of aesEncrypt_Unrolled is
  signal addroundkey0_io_s_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_s_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey0_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal nextrc0_io_ret : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal keyschedule0_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal subbytes1_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal shiftrows1_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal mixcolumns1_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey1_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal nextrc1_io_ret : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal keyschedule1_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal subbytes2_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal shiftrows2_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal mixcolumns2_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey2_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal nextrc2_io_ret : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal keyschedule2_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal subbytes3_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal shiftrows3_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal mixcolumns3_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey3_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal nextrc3_io_ret : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal keyschedule3_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal subbytes4_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal shiftrows4_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal mixcolumns4_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey4_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal nextrc4_io_ret : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal keyschedule4_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal subbytes5_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal shiftrows5_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal mixcolumns5_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey5_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal nextrc5_io_ret : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal keyschedule5_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal subbytes6_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal shiftrows6_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal mixcolumns6_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey6_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal nextrc6_io_ret : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal keyschedule6_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal subbytes7_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal shiftrows7_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal mixcolumns7_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey7_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal nextrc7_io_ret : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal keyschedule7_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal subbytes8_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal shiftrows8_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal mixcolumns8_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey8_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal nextrc8_io_ret : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal keyschedule8_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal subbytes9_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal shiftrows9_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal mixcolumns9_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey9_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal nextrc9_io_ret : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal keyschedule9_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal subbytes10_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal shiftrows10_io_ret_3_3 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_0_0 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_0_1 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_0_2 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_0_3 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_1_0 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_1_1 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_1_2 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_1_3 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_2_0 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_2_1 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_2_2 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_2_3 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_3_0 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_3_1 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_3_2 : std_logic_vector(7 downto 0);
  signal addroundkey10_io_ret_3_3 : std_logic_vector(7 downto 0);

  signal dummy : std_logic;
  signal state0_0_0 : std_logic_vector(7 downto 0);
  signal state0_0_1 : std_logic_vector(7 downto 0);
  signal state0_0_2 : std_logic_vector(7 downto 0);
  signal state0_0_3 : std_logic_vector(7 downto 0);
  signal state0_1_0 : std_logic_vector(7 downto 0);
  signal state0_1_1 : std_logic_vector(7 downto 0);
  signal state0_1_2 : std_logic_vector(7 downto 0);
  signal state0_1_3 : std_logic_vector(7 downto 0);
  signal state0_2_0 : std_logic_vector(7 downto 0);
  signal state0_2_1 : std_logic_vector(7 downto 0);
  signal state0_2_2 : std_logic_vector(7 downto 0);
  signal state0_2_3 : std_logic_vector(7 downto 0);
  signal state0_3_0 : std_logic_vector(7 downto 0);
  signal state0_3_1 : std_logic_vector(7 downto 0);
  signal state0_3_2 : std_logic_vector(7 downto 0);
  signal state0_3_3 : std_logic_vector(7 downto 0);
  signal rcs0 : std_logic_vector(7 downto 0);
  signal keys0_0_0 : std_logic_vector(7 downto 0);
  signal keys0_0_1 : std_logic_vector(7 downto 0);
  signal keys0_0_2 : std_logic_vector(7 downto 0);
  signal keys0_0_3 : std_logic_vector(7 downto 0);
  signal keys0_1_0 : std_logic_vector(7 downto 0);
  signal keys0_1_1 : std_logic_vector(7 downto 0);
  signal keys0_1_2 : std_logic_vector(7 downto 0);
  signal keys0_1_3 : std_logic_vector(7 downto 0);
  signal keys0_2_0 : std_logic_vector(7 downto 0);
  signal keys0_2_1 : std_logic_vector(7 downto 0);
  signal keys0_2_2 : std_logic_vector(7 downto 0);
  signal keys0_2_3 : std_logic_vector(7 downto 0);
  signal keys0_3_0 : std_logic_vector(7 downto 0);
  signal keys0_3_1 : std_logic_vector(7 downto 0);
  signal keys0_3_2 : std_logic_vector(7 downto 0);
  signal keys0_3_3 : std_logic_vector(7 downto 0);
  signal zz_io_ret : std_logic_vector(127 downto 0);
begin
  addroundkey0 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keys0_0_0,
      io_rk_0_1 => keys0_0_1,
      io_rk_0_2 => keys0_0_2,
      io_rk_0_3 => keys0_0_3,
      io_rk_1_0 => keys0_1_0,
      io_rk_1_1 => keys0_1_1,
      io_rk_1_2 => keys0_1_2,
      io_rk_1_3 => keys0_1_3,
      io_rk_2_0 => keys0_2_0,
      io_rk_2_1 => keys0_2_1,
      io_rk_2_2 => keys0_2_2,
      io_rk_2_3 => keys0_2_3,
      io_rk_3_0 => keys0_3_0,
      io_rk_3_1 => keys0_3_1,
      io_rk_3_2 => keys0_3_2,
      io_rk_3_3 => keys0_3_3,
      io_s_0_0 => addroundkey0_io_s_0_0,
      io_s_0_1 => addroundkey0_io_s_0_1,
      io_s_0_2 => addroundkey0_io_s_0_2,
      io_s_0_3 => addroundkey0_io_s_0_3,
      io_s_1_0 => addroundkey0_io_s_1_0,
      io_s_1_1 => addroundkey0_io_s_1_1,
      io_s_1_2 => addroundkey0_io_s_1_2,
      io_s_1_3 => addroundkey0_io_s_1_3,
      io_s_2_0 => addroundkey0_io_s_2_0,
      io_s_2_1 => addroundkey0_io_s_2_1,
      io_s_2_2 => addroundkey0_io_s_2_2,
      io_s_2_3 => addroundkey0_io_s_2_3,
      io_s_3_0 => addroundkey0_io_s_3_0,
      io_s_3_1 => addroundkey0_io_s_3_1,
      io_s_3_2 => addroundkey0_io_s_3_2,
      io_s_3_3 => addroundkey0_io_s_3_3,
      io_ret_0_0 => addroundkey0_io_ret_0_0,
      io_ret_0_1 => addroundkey0_io_ret_0_1,
      io_ret_0_2 => addroundkey0_io_ret_0_2,
      io_ret_0_3 => addroundkey0_io_ret_0_3,
      io_ret_1_0 => addroundkey0_io_ret_1_0,
      io_ret_1_1 => addroundkey0_io_ret_1_1,
      io_ret_1_2 => addroundkey0_io_ret_1_2,
      io_ret_1_3 => addroundkey0_io_ret_1_3,
      io_ret_2_0 => addroundkey0_io_ret_2_0,
      io_ret_2_1 => addroundkey0_io_ret_2_1,
      io_ret_2_2 => addroundkey0_io_ret_2_2,
      io_ret_2_3 => addroundkey0_io_ret_2_3,
      io_ret_3_0 => addroundkey0_io_ret_3_0,
      io_ret_3_1 => addroundkey0_io_ret_3_1,
      io_ret_3_2 => addroundkey0_io_ret_3_2,
      io_ret_3_3 => addroundkey0_io_ret_3_3 
    );
  nextrc0 : entity work.NextRC
    port map ( 
      io_rc => rcs0,
      io_ret => nextrc0_io_ret 
    );
  keyschedule0 : entity work.KeySchedule
    port map ( 
      io_key_0_0 => keys0_0_0,
      io_key_0_1 => keys0_0_1,
      io_key_0_2 => keys0_0_2,
      io_key_0_3 => keys0_0_3,
      io_key_1_0 => keys0_1_0,
      io_key_1_1 => keys0_1_1,
      io_key_1_2 => keys0_1_2,
      io_key_1_3 => keys0_1_3,
      io_key_2_0 => keys0_2_0,
      io_key_2_1 => keys0_2_1,
      io_key_2_2 => keys0_2_2,
      io_key_2_3 => keys0_2_3,
      io_key_3_0 => keys0_3_0,
      io_key_3_1 => keys0_3_1,
      io_key_3_2 => keys0_3_2,
      io_key_3_3 => keys0_3_3,
      io_c => rcs0,
      io_ret_0_0 => keyschedule0_io_ret_0_0,
      io_ret_0_1 => keyschedule0_io_ret_0_1,
      io_ret_0_2 => keyschedule0_io_ret_0_2,
      io_ret_0_3 => keyschedule0_io_ret_0_3,
      io_ret_1_0 => keyschedule0_io_ret_1_0,
      io_ret_1_1 => keyschedule0_io_ret_1_1,
      io_ret_1_2 => keyschedule0_io_ret_1_2,
      io_ret_1_3 => keyschedule0_io_ret_1_3,
      io_ret_2_0 => keyschedule0_io_ret_2_0,
      io_ret_2_1 => keyschedule0_io_ret_2_1,
      io_ret_2_2 => keyschedule0_io_ret_2_2,
      io_ret_2_3 => keyschedule0_io_ret_2_3,
      io_ret_3_0 => keyschedule0_io_ret_3_0,
      io_ret_3_1 => keyschedule0_io_ret_3_1,
      io_ret_3_2 => keyschedule0_io_ret_3_2,
      io_ret_3_3 => keyschedule0_io_ret_3_3 
    );
  subbytes1 : entity work.SubBytes
    port map ( 
      io_state_0_0 => state0_0_0,
      io_state_0_1 => state0_0_1,
      io_state_0_2 => state0_0_2,
      io_state_0_3 => state0_0_3,
      io_state_1_0 => state0_1_0,
      io_state_1_1 => state0_1_1,
      io_state_1_2 => state0_1_2,
      io_state_1_3 => state0_1_3,
      io_state_2_0 => state0_2_0,
      io_state_2_1 => state0_2_1,
      io_state_2_2 => state0_2_2,
      io_state_2_3 => state0_2_3,
      io_state_3_0 => state0_3_0,
      io_state_3_1 => state0_3_1,
      io_state_3_2 => state0_3_2,
      io_state_3_3 => state0_3_3,
      io_ret_0_0 => subbytes1_io_ret_0_0,
      io_ret_0_1 => subbytes1_io_ret_0_1,
      io_ret_0_2 => subbytes1_io_ret_0_2,
      io_ret_0_3 => subbytes1_io_ret_0_3,
      io_ret_1_0 => subbytes1_io_ret_1_0,
      io_ret_1_1 => subbytes1_io_ret_1_1,
      io_ret_1_2 => subbytes1_io_ret_1_2,
      io_ret_1_3 => subbytes1_io_ret_1_3,
      io_ret_2_0 => subbytes1_io_ret_2_0,
      io_ret_2_1 => subbytes1_io_ret_2_1,
      io_ret_2_2 => subbytes1_io_ret_2_2,
      io_ret_2_3 => subbytes1_io_ret_2_3,
      io_ret_3_0 => subbytes1_io_ret_3_0,
      io_ret_3_1 => subbytes1_io_ret_3_1,
      io_ret_3_2 => subbytes1_io_ret_3_2,
      io_ret_3_3 => subbytes1_io_ret_3_3 
    );
  shiftrows1 : entity work.ShiftRows
    port map ( 
      io_state_0_0 => subbytes1_io_ret_0_0,
      io_state_0_1 => subbytes1_io_ret_0_1,
      io_state_0_2 => subbytes1_io_ret_0_2,
      io_state_0_3 => subbytes1_io_ret_0_3,
      io_state_1_0 => subbytes1_io_ret_1_0,
      io_state_1_1 => subbytes1_io_ret_1_1,
      io_state_1_2 => subbytes1_io_ret_1_2,
      io_state_1_3 => subbytes1_io_ret_1_3,
      io_state_2_0 => subbytes1_io_ret_2_0,
      io_state_2_1 => subbytes1_io_ret_2_1,
      io_state_2_2 => subbytes1_io_ret_2_2,
      io_state_2_3 => subbytes1_io_ret_2_3,
      io_state_3_0 => subbytes1_io_ret_3_0,
      io_state_3_1 => subbytes1_io_ret_3_1,
      io_state_3_2 => subbytes1_io_ret_3_2,
      io_state_3_3 => subbytes1_io_ret_3_3,
      io_ret_0_0 => shiftrows1_io_ret_0_0,
      io_ret_0_1 => shiftrows1_io_ret_0_1,
      io_ret_0_2 => shiftrows1_io_ret_0_2,
      io_ret_0_3 => shiftrows1_io_ret_0_3,
      io_ret_1_0 => shiftrows1_io_ret_1_0,
      io_ret_1_1 => shiftrows1_io_ret_1_1,
      io_ret_1_2 => shiftrows1_io_ret_1_2,
      io_ret_1_3 => shiftrows1_io_ret_1_3,
      io_ret_2_0 => shiftrows1_io_ret_2_0,
      io_ret_2_1 => shiftrows1_io_ret_2_1,
      io_ret_2_2 => shiftrows1_io_ret_2_2,
      io_ret_2_3 => shiftrows1_io_ret_2_3,
      io_ret_3_0 => shiftrows1_io_ret_3_0,
      io_ret_3_1 => shiftrows1_io_ret_3_1,
      io_ret_3_2 => shiftrows1_io_ret_3_2,
      io_ret_3_3 => shiftrows1_io_ret_3_3 
    );
  mixcolumns1 : entity work.MixColumns
    port map ( 
      io_state_0_0 => shiftrows1_io_ret_0_0,
      io_state_0_1 => shiftrows1_io_ret_0_1,
      io_state_0_2 => shiftrows1_io_ret_0_2,
      io_state_0_3 => shiftrows1_io_ret_0_3,
      io_state_1_0 => shiftrows1_io_ret_1_0,
      io_state_1_1 => shiftrows1_io_ret_1_1,
      io_state_1_2 => shiftrows1_io_ret_1_2,
      io_state_1_3 => shiftrows1_io_ret_1_3,
      io_state_2_0 => shiftrows1_io_ret_2_0,
      io_state_2_1 => shiftrows1_io_ret_2_1,
      io_state_2_2 => shiftrows1_io_ret_2_2,
      io_state_2_3 => shiftrows1_io_ret_2_3,
      io_state_3_0 => shiftrows1_io_ret_3_0,
      io_state_3_1 => shiftrows1_io_ret_3_1,
      io_state_3_2 => shiftrows1_io_ret_3_2,
      io_state_3_3 => shiftrows1_io_ret_3_3,
      io_ret_0_0 => mixcolumns1_io_ret_0_0,
      io_ret_0_1 => mixcolumns1_io_ret_0_1,
      io_ret_0_2 => mixcolumns1_io_ret_0_2,
      io_ret_0_3 => mixcolumns1_io_ret_0_3,
      io_ret_1_0 => mixcolumns1_io_ret_1_0,
      io_ret_1_1 => mixcolumns1_io_ret_1_1,
      io_ret_1_2 => mixcolumns1_io_ret_1_2,
      io_ret_1_3 => mixcolumns1_io_ret_1_3,
      io_ret_2_0 => mixcolumns1_io_ret_2_0,
      io_ret_2_1 => mixcolumns1_io_ret_2_1,
      io_ret_2_2 => mixcolumns1_io_ret_2_2,
      io_ret_2_3 => mixcolumns1_io_ret_2_3,
      io_ret_3_0 => mixcolumns1_io_ret_3_0,
      io_ret_3_1 => mixcolumns1_io_ret_3_1,
      io_ret_3_2 => mixcolumns1_io_ret_3_2,
      io_ret_3_3 => mixcolumns1_io_ret_3_3 
    );
  addroundkey1 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keyschedule0_io_ret_0_0,
      io_rk_0_1 => keyschedule0_io_ret_0_1,
      io_rk_0_2 => keyschedule0_io_ret_0_2,
      io_rk_0_3 => keyschedule0_io_ret_0_3,
      io_rk_1_0 => keyschedule0_io_ret_1_0,
      io_rk_1_1 => keyschedule0_io_ret_1_1,
      io_rk_1_2 => keyschedule0_io_ret_1_2,
      io_rk_1_3 => keyschedule0_io_ret_1_3,
      io_rk_2_0 => keyschedule0_io_ret_2_0,
      io_rk_2_1 => keyschedule0_io_ret_2_1,
      io_rk_2_2 => keyschedule0_io_ret_2_2,
      io_rk_2_3 => keyschedule0_io_ret_2_3,
      io_rk_3_0 => keyschedule0_io_ret_3_0,
      io_rk_3_1 => keyschedule0_io_ret_3_1,
      io_rk_3_2 => keyschedule0_io_ret_3_2,
      io_rk_3_3 => keyschedule0_io_ret_3_3,
      io_s_0_0 => mixcolumns1_io_ret_0_0,
      io_s_0_1 => mixcolumns1_io_ret_0_1,
      io_s_0_2 => mixcolumns1_io_ret_0_2,
      io_s_0_3 => mixcolumns1_io_ret_0_3,
      io_s_1_0 => mixcolumns1_io_ret_1_0,
      io_s_1_1 => mixcolumns1_io_ret_1_1,
      io_s_1_2 => mixcolumns1_io_ret_1_2,
      io_s_1_3 => mixcolumns1_io_ret_1_3,
      io_s_2_0 => mixcolumns1_io_ret_2_0,
      io_s_2_1 => mixcolumns1_io_ret_2_1,
      io_s_2_2 => mixcolumns1_io_ret_2_2,
      io_s_2_3 => mixcolumns1_io_ret_2_3,
      io_s_3_0 => mixcolumns1_io_ret_3_0,
      io_s_3_1 => mixcolumns1_io_ret_3_1,
      io_s_3_2 => mixcolumns1_io_ret_3_2,
      io_s_3_3 => mixcolumns1_io_ret_3_3,
      io_ret_0_0 => addroundkey1_io_ret_0_0,
      io_ret_0_1 => addroundkey1_io_ret_0_1,
      io_ret_0_2 => addroundkey1_io_ret_0_2,
      io_ret_0_3 => addroundkey1_io_ret_0_3,
      io_ret_1_0 => addroundkey1_io_ret_1_0,
      io_ret_1_1 => addroundkey1_io_ret_1_1,
      io_ret_1_2 => addroundkey1_io_ret_1_2,
      io_ret_1_3 => addroundkey1_io_ret_1_3,
      io_ret_2_0 => addroundkey1_io_ret_2_0,
      io_ret_2_1 => addroundkey1_io_ret_2_1,
      io_ret_2_2 => addroundkey1_io_ret_2_2,
      io_ret_2_3 => addroundkey1_io_ret_2_3,
      io_ret_3_0 => addroundkey1_io_ret_3_0,
      io_ret_3_1 => addroundkey1_io_ret_3_1,
      io_ret_3_2 => addroundkey1_io_ret_3_2,
      io_ret_3_3 => addroundkey1_io_ret_3_3 
    );
  nextrc1 : entity work.NextRC
    port map ( 
      io_rc => nextrc0_io_ret,
      io_ret => nextrc1_io_ret 
    );
  keyschedule1 : entity work.KeySchedule
    port map ( 
      io_key_0_0 => keyschedule0_io_ret_0_0,
      io_key_0_1 => keyschedule0_io_ret_0_1,
      io_key_0_2 => keyschedule0_io_ret_0_2,
      io_key_0_3 => keyschedule0_io_ret_0_3,
      io_key_1_0 => keyschedule0_io_ret_1_0,
      io_key_1_1 => keyschedule0_io_ret_1_1,
      io_key_1_2 => keyschedule0_io_ret_1_2,
      io_key_1_3 => keyschedule0_io_ret_1_3,
      io_key_2_0 => keyschedule0_io_ret_2_0,
      io_key_2_1 => keyschedule0_io_ret_2_1,
      io_key_2_2 => keyschedule0_io_ret_2_2,
      io_key_2_3 => keyschedule0_io_ret_2_3,
      io_key_3_0 => keyschedule0_io_ret_3_0,
      io_key_3_1 => keyschedule0_io_ret_3_1,
      io_key_3_2 => keyschedule0_io_ret_3_2,
      io_key_3_3 => keyschedule0_io_ret_3_3,
      io_c => nextrc0_io_ret,
      io_ret_0_0 => keyschedule1_io_ret_0_0,
      io_ret_0_1 => keyschedule1_io_ret_0_1,
      io_ret_0_2 => keyschedule1_io_ret_0_2,
      io_ret_0_3 => keyschedule1_io_ret_0_3,
      io_ret_1_0 => keyschedule1_io_ret_1_0,
      io_ret_1_1 => keyschedule1_io_ret_1_1,
      io_ret_1_2 => keyschedule1_io_ret_1_2,
      io_ret_1_3 => keyschedule1_io_ret_1_3,
      io_ret_2_0 => keyschedule1_io_ret_2_0,
      io_ret_2_1 => keyschedule1_io_ret_2_1,
      io_ret_2_2 => keyschedule1_io_ret_2_2,
      io_ret_2_3 => keyschedule1_io_ret_2_3,
      io_ret_3_0 => keyschedule1_io_ret_3_0,
      io_ret_3_1 => keyschedule1_io_ret_3_1,
      io_ret_3_2 => keyschedule1_io_ret_3_2,
      io_ret_3_3 => keyschedule1_io_ret_3_3 
    );
  subbytes2 : entity work.SubBytes
    port map ( 
      io_state_0_0 => addroundkey1_io_ret_0_0,
      io_state_0_1 => addroundkey1_io_ret_0_1,
      io_state_0_2 => addroundkey1_io_ret_0_2,
      io_state_0_3 => addroundkey1_io_ret_0_3,
      io_state_1_0 => addroundkey1_io_ret_1_0,
      io_state_1_1 => addroundkey1_io_ret_1_1,
      io_state_1_2 => addroundkey1_io_ret_1_2,
      io_state_1_3 => addroundkey1_io_ret_1_3,
      io_state_2_0 => addroundkey1_io_ret_2_0,
      io_state_2_1 => addroundkey1_io_ret_2_1,
      io_state_2_2 => addroundkey1_io_ret_2_2,
      io_state_2_3 => addroundkey1_io_ret_2_3,
      io_state_3_0 => addroundkey1_io_ret_3_0,
      io_state_3_1 => addroundkey1_io_ret_3_1,
      io_state_3_2 => addroundkey1_io_ret_3_2,
      io_state_3_3 => addroundkey1_io_ret_3_3,
      io_ret_0_0 => subbytes2_io_ret_0_0,
      io_ret_0_1 => subbytes2_io_ret_0_1,
      io_ret_0_2 => subbytes2_io_ret_0_2,
      io_ret_0_3 => subbytes2_io_ret_0_3,
      io_ret_1_0 => subbytes2_io_ret_1_0,
      io_ret_1_1 => subbytes2_io_ret_1_1,
      io_ret_1_2 => subbytes2_io_ret_1_2,
      io_ret_1_3 => subbytes2_io_ret_1_3,
      io_ret_2_0 => subbytes2_io_ret_2_0,
      io_ret_2_1 => subbytes2_io_ret_2_1,
      io_ret_2_2 => subbytes2_io_ret_2_2,
      io_ret_2_3 => subbytes2_io_ret_2_3,
      io_ret_3_0 => subbytes2_io_ret_3_0,
      io_ret_3_1 => subbytes2_io_ret_3_1,
      io_ret_3_2 => subbytes2_io_ret_3_2,
      io_ret_3_3 => subbytes2_io_ret_3_3 
    );
  shiftrows2 : entity work.ShiftRows
    port map ( 
      io_state_0_0 => subbytes2_io_ret_0_0,
      io_state_0_1 => subbytes2_io_ret_0_1,
      io_state_0_2 => subbytes2_io_ret_0_2,
      io_state_0_3 => subbytes2_io_ret_0_3,
      io_state_1_0 => subbytes2_io_ret_1_0,
      io_state_1_1 => subbytes2_io_ret_1_1,
      io_state_1_2 => subbytes2_io_ret_1_2,
      io_state_1_3 => subbytes2_io_ret_1_3,
      io_state_2_0 => subbytes2_io_ret_2_0,
      io_state_2_1 => subbytes2_io_ret_2_1,
      io_state_2_2 => subbytes2_io_ret_2_2,
      io_state_2_3 => subbytes2_io_ret_2_3,
      io_state_3_0 => subbytes2_io_ret_3_0,
      io_state_3_1 => subbytes2_io_ret_3_1,
      io_state_3_2 => subbytes2_io_ret_3_2,
      io_state_3_3 => subbytes2_io_ret_3_3,
      io_ret_0_0 => shiftrows2_io_ret_0_0,
      io_ret_0_1 => shiftrows2_io_ret_0_1,
      io_ret_0_2 => shiftrows2_io_ret_0_2,
      io_ret_0_3 => shiftrows2_io_ret_0_3,
      io_ret_1_0 => shiftrows2_io_ret_1_0,
      io_ret_1_1 => shiftrows2_io_ret_1_1,
      io_ret_1_2 => shiftrows2_io_ret_1_2,
      io_ret_1_3 => shiftrows2_io_ret_1_3,
      io_ret_2_0 => shiftrows2_io_ret_2_0,
      io_ret_2_1 => shiftrows2_io_ret_2_1,
      io_ret_2_2 => shiftrows2_io_ret_2_2,
      io_ret_2_3 => shiftrows2_io_ret_2_3,
      io_ret_3_0 => shiftrows2_io_ret_3_0,
      io_ret_3_1 => shiftrows2_io_ret_3_1,
      io_ret_3_2 => shiftrows2_io_ret_3_2,
      io_ret_3_3 => shiftrows2_io_ret_3_3 
    );
  mixcolumns2 : entity work.MixColumns
    port map ( 
      io_state_0_0 => shiftrows2_io_ret_0_0,
      io_state_0_1 => shiftrows2_io_ret_0_1,
      io_state_0_2 => shiftrows2_io_ret_0_2,
      io_state_0_3 => shiftrows2_io_ret_0_3,
      io_state_1_0 => shiftrows2_io_ret_1_0,
      io_state_1_1 => shiftrows2_io_ret_1_1,
      io_state_1_2 => shiftrows2_io_ret_1_2,
      io_state_1_3 => shiftrows2_io_ret_1_3,
      io_state_2_0 => shiftrows2_io_ret_2_0,
      io_state_2_1 => shiftrows2_io_ret_2_1,
      io_state_2_2 => shiftrows2_io_ret_2_2,
      io_state_2_3 => shiftrows2_io_ret_2_3,
      io_state_3_0 => shiftrows2_io_ret_3_0,
      io_state_3_1 => shiftrows2_io_ret_3_1,
      io_state_3_2 => shiftrows2_io_ret_3_2,
      io_state_3_3 => shiftrows2_io_ret_3_3,
      io_ret_0_0 => mixcolumns2_io_ret_0_0,
      io_ret_0_1 => mixcolumns2_io_ret_0_1,
      io_ret_0_2 => mixcolumns2_io_ret_0_2,
      io_ret_0_3 => mixcolumns2_io_ret_0_3,
      io_ret_1_0 => mixcolumns2_io_ret_1_0,
      io_ret_1_1 => mixcolumns2_io_ret_1_1,
      io_ret_1_2 => mixcolumns2_io_ret_1_2,
      io_ret_1_3 => mixcolumns2_io_ret_1_3,
      io_ret_2_0 => mixcolumns2_io_ret_2_0,
      io_ret_2_1 => mixcolumns2_io_ret_2_1,
      io_ret_2_2 => mixcolumns2_io_ret_2_2,
      io_ret_2_3 => mixcolumns2_io_ret_2_3,
      io_ret_3_0 => mixcolumns2_io_ret_3_0,
      io_ret_3_1 => mixcolumns2_io_ret_3_1,
      io_ret_3_2 => mixcolumns2_io_ret_3_2,
      io_ret_3_3 => mixcolumns2_io_ret_3_3 
    );
  addroundkey2 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keyschedule1_io_ret_0_0,
      io_rk_0_1 => keyschedule1_io_ret_0_1,
      io_rk_0_2 => keyschedule1_io_ret_0_2,
      io_rk_0_3 => keyschedule1_io_ret_0_3,
      io_rk_1_0 => keyschedule1_io_ret_1_0,
      io_rk_1_1 => keyschedule1_io_ret_1_1,
      io_rk_1_2 => keyschedule1_io_ret_1_2,
      io_rk_1_3 => keyschedule1_io_ret_1_3,
      io_rk_2_0 => keyschedule1_io_ret_2_0,
      io_rk_2_1 => keyschedule1_io_ret_2_1,
      io_rk_2_2 => keyschedule1_io_ret_2_2,
      io_rk_2_3 => keyschedule1_io_ret_2_3,
      io_rk_3_0 => keyschedule1_io_ret_3_0,
      io_rk_3_1 => keyschedule1_io_ret_3_1,
      io_rk_3_2 => keyschedule1_io_ret_3_2,
      io_rk_3_3 => keyschedule1_io_ret_3_3,
      io_s_0_0 => mixcolumns2_io_ret_0_0,
      io_s_0_1 => mixcolumns2_io_ret_0_1,
      io_s_0_2 => mixcolumns2_io_ret_0_2,
      io_s_0_3 => mixcolumns2_io_ret_0_3,
      io_s_1_0 => mixcolumns2_io_ret_1_0,
      io_s_1_1 => mixcolumns2_io_ret_1_1,
      io_s_1_2 => mixcolumns2_io_ret_1_2,
      io_s_1_3 => mixcolumns2_io_ret_1_3,
      io_s_2_0 => mixcolumns2_io_ret_2_0,
      io_s_2_1 => mixcolumns2_io_ret_2_1,
      io_s_2_2 => mixcolumns2_io_ret_2_2,
      io_s_2_3 => mixcolumns2_io_ret_2_3,
      io_s_3_0 => mixcolumns2_io_ret_3_0,
      io_s_3_1 => mixcolumns2_io_ret_3_1,
      io_s_3_2 => mixcolumns2_io_ret_3_2,
      io_s_3_3 => mixcolumns2_io_ret_3_3,
      io_ret_0_0 => addroundkey2_io_ret_0_0,
      io_ret_0_1 => addroundkey2_io_ret_0_1,
      io_ret_0_2 => addroundkey2_io_ret_0_2,
      io_ret_0_3 => addroundkey2_io_ret_0_3,
      io_ret_1_0 => addroundkey2_io_ret_1_0,
      io_ret_1_1 => addroundkey2_io_ret_1_1,
      io_ret_1_2 => addroundkey2_io_ret_1_2,
      io_ret_1_3 => addroundkey2_io_ret_1_3,
      io_ret_2_0 => addroundkey2_io_ret_2_0,
      io_ret_2_1 => addroundkey2_io_ret_2_1,
      io_ret_2_2 => addroundkey2_io_ret_2_2,
      io_ret_2_3 => addroundkey2_io_ret_2_3,
      io_ret_3_0 => addroundkey2_io_ret_3_0,
      io_ret_3_1 => addroundkey2_io_ret_3_1,
      io_ret_3_2 => addroundkey2_io_ret_3_2,
      io_ret_3_3 => addroundkey2_io_ret_3_3 
    );
  nextrc2 : entity work.NextRC
    port map ( 
      io_rc => nextrc1_io_ret,
      io_ret => nextrc2_io_ret 
    );
  keyschedule2 : entity work.KeySchedule
    port map ( 
      io_key_0_0 => keyschedule1_io_ret_0_0,
      io_key_0_1 => keyschedule1_io_ret_0_1,
      io_key_0_2 => keyschedule1_io_ret_0_2,
      io_key_0_3 => keyschedule1_io_ret_0_3,
      io_key_1_0 => keyschedule1_io_ret_1_0,
      io_key_1_1 => keyschedule1_io_ret_1_1,
      io_key_1_2 => keyschedule1_io_ret_1_2,
      io_key_1_3 => keyschedule1_io_ret_1_3,
      io_key_2_0 => keyschedule1_io_ret_2_0,
      io_key_2_1 => keyschedule1_io_ret_2_1,
      io_key_2_2 => keyschedule1_io_ret_2_2,
      io_key_2_3 => keyschedule1_io_ret_2_3,
      io_key_3_0 => keyschedule1_io_ret_3_0,
      io_key_3_1 => keyschedule1_io_ret_3_1,
      io_key_3_2 => keyschedule1_io_ret_3_2,
      io_key_3_3 => keyschedule1_io_ret_3_3,
      io_c => nextrc1_io_ret,
      io_ret_0_0 => keyschedule2_io_ret_0_0,
      io_ret_0_1 => keyschedule2_io_ret_0_1,
      io_ret_0_2 => keyschedule2_io_ret_0_2,
      io_ret_0_3 => keyschedule2_io_ret_0_3,
      io_ret_1_0 => keyschedule2_io_ret_1_0,
      io_ret_1_1 => keyschedule2_io_ret_1_1,
      io_ret_1_2 => keyschedule2_io_ret_1_2,
      io_ret_1_3 => keyschedule2_io_ret_1_3,
      io_ret_2_0 => keyschedule2_io_ret_2_0,
      io_ret_2_1 => keyschedule2_io_ret_2_1,
      io_ret_2_2 => keyschedule2_io_ret_2_2,
      io_ret_2_3 => keyschedule2_io_ret_2_3,
      io_ret_3_0 => keyschedule2_io_ret_3_0,
      io_ret_3_1 => keyschedule2_io_ret_3_1,
      io_ret_3_2 => keyschedule2_io_ret_3_2,
      io_ret_3_3 => keyschedule2_io_ret_3_3 
    );
  subbytes3 : entity work.SubBytes
    port map ( 
      io_state_0_0 => addroundkey2_io_ret_0_0,
      io_state_0_1 => addroundkey2_io_ret_0_1,
      io_state_0_2 => addroundkey2_io_ret_0_2,
      io_state_0_3 => addroundkey2_io_ret_0_3,
      io_state_1_0 => addroundkey2_io_ret_1_0,
      io_state_1_1 => addroundkey2_io_ret_1_1,
      io_state_1_2 => addroundkey2_io_ret_1_2,
      io_state_1_3 => addroundkey2_io_ret_1_3,
      io_state_2_0 => addroundkey2_io_ret_2_0,
      io_state_2_1 => addroundkey2_io_ret_2_1,
      io_state_2_2 => addroundkey2_io_ret_2_2,
      io_state_2_3 => addroundkey2_io_ret_2_3,
      io_state_3_0 => addroundkey2_io_ret_3_0,
      io_state_3_1 => addroundkey2_io_ret_3_1,
      io_state_3_2 => addroundkey2_io_ret_3_2,
      io_state_3_3 => addroundkey2_io_ret_3_3,
      io_ret_0_0 => subbytes3_io_ret_0_0,
      io_ret_0_1 => subbytes3_io_ret_0_1,
      io_ret_0_2 => subbytes3_io_ret_0_2,
      io_ret_0_3 => subbytes3_io_ret_0_3,
      io_ret_1_0 => subbytes3_io_ret_1_0,
      io_ret_1_1 => subbytes3_io_ret_1_1,
      io_ret_1_2 => subbytes3_io_ret_1_2,
      io_ret_1_3 => subbytes3_io_ret_1_3,
      io_ret_2_0 => subbytes3_io_ret_2_0,
      io_ret_2_1 => subbytes3_io_ret_2_1,
      io_ret_2_2 => subbytes3_io_ret_2_2,
      io_ret_2_3 => subbytes3_io_ret_2_3,
      io_ret_3_0 => subbytes3_io_ret_3_0,
      io_ret_3_1 => subbytes3_io_ret_3_1,
      io_ret_3_2 => subbytes3_io_ret_3_2,
      io_ret_3_3 => subbytes3_io_ret_3_3 
    );
  shiftrows3 : entity work.ShiftRows
    port map ( 
      io_state_0_0 => subbytes3_io_ret_0_0,
      io_state_0_1 => subbytes3_io_ret_0_1,
      io_state_0_2 => subbytes3_io_ret_0_2,
      io_state_0_3 => subbytes3_io_ret_0_3,
      io_state_1_0 => subbytes3_io_ret_1_0,
      io_state_1_1 => subbytes3_io_ret_1_1,
      io_state_1_2 => subbytes3_io_ret_1_2,
      io_state_1_3 => subbytes3_io_ret_1_3,
      io_state_2_0 => subbytes3_io_ret_2_0,
      io_state_2_1 => subbytes3_io_ret_2_1,
      io_state_2_2 => subbytes3_io_ret_2_2,
      io_state_2_3 => subbytes3_io_ret_2_3,
      io_state_3_0 => subbytes3_io_ret_3_0,
      io_state_3_1 => subbytes3_io_ret_3_1,
      io_state_3_2 => subbytes3_io_ret_3_2,
      io_state_3_3 => subbytes3_io_ret_3_3,
      io_ret_0_0 => shiftrows3_io_ret_0_0,
      io_ret_0_1 => shiftrows3_io_ret_0_1,
      io_ret_0_2 => shiftrows3_io_ret_0_2,
      io_ret_0_3 => shiftrows3_io_ret_0_3,
      io_ret_1_0 => shiftrows3_io_ret_1_0,
      io_ret_1_1 => shiftrows3_io_ret_1_1,
      io_ret_1_2 => shiftrows3_io_ret_1_2,
      io_ret_1_3 => shiftrows3_io_ret_1_3,
      io_ret_2_0 => shiftrows3_io_ret_2_0,
      io_ret_2_1 => shiftrows3_io_ret_2_1,
      io_ret_2_2 => shiftrows3_io_ret_2_2,
      io_ret_2_3 => shiftrows3_io_ret_2_3,
      io_ret_3_0 => shiftrows3_io_ret_3_0,
      io_ret_3_1 => shiftrows3_io_ret_3_1,
      io_ret_3_2 => shiftrows3_io_ret_3_2,
      io_ret_3_3 => shiftrows3_io_ret_3_3 
    );
  mixcolumns3 : entity work.MixColumns
    port map ( 
      io_state_0_0 => shiftrows3_io_ret_0_0,
      io_state_0_1 => shiftrows3_io_ret_0_1,
      io_state_0_2 => shiftrows3_io_ret_0_2,
      io_state_0_3 => shiftrows3_io_ret_0_3,
      io_state_1_0 => shiftrows3_io_ret_1_0,
      io_state_1_1 => shiftrows3_io_ret_1_1,
      io_state_1_2 => shiftrows3_io_ret_1_2,
      io_state_1_3 => shiftrows3_io_ret_1_3,
      io_state_2_0 => shiftrows3_io_ret_2_0,
      io_state_2_1 => shiftrows3_io_ret_2_1,
      io_state_2_2 => shiftrows3_io_ret_2_2,
      io_state_2_3 => shiftrows3_io_ret_2_3,
      io_state_3_0 => shiftrows3_io_ret_3_0,
      io_state_3_1 => shiftrows3_io_ret_3_1,
      io_state_3_2 => shiftrows3_io_ret_3_2,
      io_state_3_3 => shiftrows3_io_ret_3_3,
      io_ret_0_0 => mixcolumns3_io_ret_0_0,
      io_ret_0_1 => mixcolumns3_io_ret_0_1,
      io_ret_0_2 => mixcolumns3_io_ret_0_2,
      io_ret_0_3 => mixcolumns3_io_ret_0_3,
      io_ret_1_0 => mixcolumns3_io_ret_1_0,
      io_ret_1_1 => mixcolumns3_io_ret_1_1,
      io_ret_1_2 => mixcolumns3_io_ret_1_2,
      io_ret_1_3 => mixcolumns3_io_ret_1_3,
      io_ret_2_0 => mixcolumns3_io_ret_2_0,
      io_ret_2_1 => mixcolumns3_io_ret_2_1,
      io_ret_2_2 => mixcolumns3_io_ret_2_2,
      io_ret_2_3 => mixcolumns3_io_ret_2_3,
      io_ret_3_0 => mixcolumns3_io_ret_3_0,
      io_ret_3_1 => mixcolumns3_io_ret_3_1,
      io_ret_3_2 => mixcolumns3_io_ret_3_2,
      io_ret_3_3 => mixcolumns3_io_ret_3_3 
    );
  addroundkey3 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keyschedule2_io_ret_0_0,
      io_rk_0_1 => keyschedule2_io_ret_0_1,
      io_rk_0_2 => keyschedule2_io_ret_0_2,
      io_rk_0_3 => keyschedule2_io_ret_0_3,
      io_rk_1_0 => keyschedule2_io_ret_1_0,
      io_rk_1_1 => keyschedule2_io_ret_1_1,
      io_rk_1_2 => keyschedule2_io_ret_1_2,
      io_rk_1_3 => keyschedule2_io_ret_1_3,
      io_rk_2_0 => keyschedule2_io_ret_2_0,
      io_rk_2_1 => keyschedule2_io_ret_2_1,
      io_rk_2_2 => keyschedule2_io_ret_2_2,
      io_rk_2_3 => keyschedule2_io_ret_2_3,
      io_rk_3_0 => keyschedule2_io_ret_3_0,
      io_rk_3_1 => keyschedule2_io_ret_3_1,
      io_rk_3_2 => keyschedule2_io_ret_3_2,
      io_rk_3_3 => keyschedule2_io_ret_3_3,
      io_s_0_0 => mixcolumns3_io_ret_0_0,
      io_s_0_1 => mixcolumns3_io_ret_0_1,
      io_s_0_2 => mixcolumns3_io_ret_0_2,
      io_s_0_3 => mixcolumns3_io_ret_0_3,
      io_s_1_0 => mixcolumns3_io_ret_1_0,
      io_s_1_1 => mixcolumns3_io_ret_1_1,
      io_s_1_2 => mixcolumns3_io_ret_1_2,
      io_s_1_3 => mixcolumns3_io_ret_1_3,
      io_s_2_0 => mixcolumns3_io_ret_2_0,
      io_s_2_1 => mixcolumns3_io_ret_2_1,
      io_s_2_2 => mixcolumns3_io_ret_2_2,
      io_s_2_3 => mixcolumns3_io_ret_2_3,
      io_s_3_0 => mixcolumns3_io_ret_3_0,
      io_s_3_1 => mixcolumns3_io_ret_3_1,
      io_s_3_2 => mixcolumns3_io_ret_3_2,
      io_s_3_3 => mixcolumns3_io_ret_3_3,
      io_ret_0_0 => addroundkey3_io_ret_0_0,
      io_ret_0_1 => addroundkey3_io_ret_0_1,
      io_ret_0_2 => addroundkey3_io_ret_0_2,
      io_ret_0_3 => addroundkey3_io_ret_0_3,
      io_ret_1_0 => addroundkey3_io_ret_1_0,
      io_ret_1_1 => addroundkey3_io_ret_1_1,
      io_ret_1_2 => addroundkey3_io_ret_1_2,
      io_ret_1_3 => addroundkey3_io_ret_1_3,
      io_ret_2_0 => addroundkey3_io_ret_2_0,
      io_ret_2_1 => addroundkey3_io_ret_2_1,
      io_ret_2_2 => addroundkey3_io_ret_2_2,
      io_ret_2_3 => addroundkey3_io_ret_2_3,
      io_ret_3_0 => addroundkey3_io_ret_3_0,
      io_ret_3_1 => addroundkey3_io_ret_3_1,
      io_ret_3_2 => addroundkey3_io_ret_3_2,
      io_ret_3_3 => addroundkey3_io_ret_3_3 
    );
  nextrc3 : entity work.NextRC
    port map ( 
      io_rc => nextrc2_io_ret,
      io_ret => nextrc3_io_ret 
    );
  keyschedule3 : entity work.KeySchedule
    port map ( 
      io_key_0_0 => keyschedule2_io_ret_0_0,
      io_key_0_1 => keyschedule2_io_ret_0_1,
      io_key_0_2 => keyschedule2_io_ret_0_2,
      io_key_0_3 => keyschedule2_io_ret_0_3,
      io_key_1_0 => keyschedule2_io_ret_1_0,
      io_key_1_1 => keyschedule2_io_ret_1_1,
      io_key_1_2 => keyschedule2_io_ret_1_2,
      io_key_1_3 => keyschedule2_io_ret_1_3,
      io_key_2_0 => keyschedule2_io_ret_2_0,
      io_key_2_1 => keyschedule2_io_ret_2_1,
      io_key_2_2 => keyschedule2_io_ret_2_2,
      io_key_2_3 => keyschedule2_io_ret_2_3,
      io_key_3_0 => keyschedule2_io_ret_3_0,
      io_key_3_1 => keyschedule2_io_ret_3_1,
      io_key_3_2 => keyschedule2_io_ret_3_2,
      io_key_3_3 => keyschedule2_io_ret_3_3,
      io_c => nextrc2_io_ret,
      io_ret_0_0 => keyschedule3_io_ret_0_0,
      io_ret_0_1 => keyschedule3_io_ret_0_1,
      io_ret_0_2 => keyschedule3_io_ret_0_2,
      io_ret_0_3 => keyschedule3_io_ret_0_3,
      io_ret_1_0 => keyschedule3_io_ret_1_0,
      io_ret_1_1 => keyschedule3_io_ret_1_1,
      io_ret_1_2 => keyschedule3_io_ret_1_2,
      io_ret_1_3 => keyschedule3_io_ret_1_3,
      io_ret_2_0 => keyschedule3_io_ret_2_0,
      io_ret_2_1 => keyschedule3_io_ret_2_1,
      io_ret_2_2 => keyschedule3_io_ret_2_2,
      io_ret_2_3 => keyschedule3_io_ret_2_3,
      io_ret_3_0 => keyschedule3_io_ret_3_0,
      io_ret_3_1 => keyschedule3_io_ret_3_1,
      io_ret_3_2 => keyschedule3_io_ret_3_2,
      io_ret_3_3 => keyschedule3_io_ret_3_3 
    );
  subbytes4 : entity work.SubBytes
    port map ( 
      io_state_0_0 => addroundkey3_io_ret_0_0,
      io_state_0_1 => addroundkey3_io_ret_0_1,
      io_state_0_2 => addroundkey3_io_ret_0_2,
      io_state_0_3 => addroundkey3_io_ret_0_3,
      io_state_1_0 => addroundkey3_io_ret_1_0,
      io_state_1_1 => addroundkey3_io_ret_1_1,
      io_state_1_2 => addroundkey3_io_ret_1_2,
      io_state_1_3 => addroundkey3_io_ret_1_3,
      io_state_2_0 => addroundkey3_io_ret_2_0,
      io_state_2_1 => addroundkey3_io_ret_2_1,
      io_state_2_2 => addroundkey3_io_ret_2_2,
      io_state_2_3 => addroundkey3_io_ret_2_3,
      io_state_3_0 => addroundkey3_io_ret_3_0,
      io_state_3_1 => addroundkey3_io_ret_3_1,
      io_state_3_2 => addroundkey3_io_ret_3_2,
      io_state_3_3 => addroundkey3_io_ret_3_3,
      io_ret_0_0 => subbytes4_io_ret_0_0,
      io_ret_0_1 => subbytes4_io_ret_0_1,
      io_ret_0_2 => subbytes4_io_ret_0_2,
      io_ret_0_3 => subbytes4_io_ret_0_3,
      io_ret_1_0 => subbytes4_io_ret_1_0,
      io_ret_1_1 => subbytes4_io_ret_1_1,
      io_ret_1_2 => subbytes4_io_ret_1_2,
      io_ret_1_3 => subbytes4_io_ret_1_3,
      io_ret_2_0 => subbytes4_io_ret_2_0,
      io_ret_2_1 => subbytes4_io_ret_2_1,
      io_ret_2_2 => subbytes4_io_ret_2_2,
      io_ret_2_3 => subbytes4_io_ret_2_3,
      io_ret_3_0 => subbytes4_io_ret_3_0,
      io_ret_3_1 => subbytes4_io_ret_3_1,
      io_ret_3_2 => subbytes4_io_ret_3_2,
      io_ret_3_3 => subbytes4_io_ret_3_3 
    );
  shiftrows4 : entity work.ShiftRows
    port map ( 
      io_state_0_0 => subbytes4_io_ret_0_0,
      io_state_0_1 => subbytes4_io_ret_0_1,
      io_state_0_2 => subbytes4_io_ret_0_2,
      io_state_0_3 => subbytes4_io_ret_0_3,
      io_state_1_0 => subbytes4_io_ret_1_0,
      io_state_1_1 => subbytes4_io_ret_1_1,
      io_state_1_2 => subbytes4_io_ret_1_2,
      io_state_1_3 => subbytes4_io_ret_1_3,
      io_state_2_0 => subbytes4_io_ret_2_0,
      io_state_2_1 => subbytes4_io_ret_2_1,
      io_state_2_2 => subbytes4_io_ret_2_2,
      io_state_2_3 => subbytes4_io_ret_2_3,
      io_state_3_0 => subbytes4_io_ret_3_0,
      io_state_3_1 => subbytes4_io_ret_3_1,
      io_state_3_2 => subbytes4_io_ret_3_2,
      io_state_3_3 => subbytes4_io_ret_3_3,
      io_ret_0_0 => shiftrows4_io_ret_0_0,
      io_ret_0_1 => shiftrows4_io_ret_0_1,
      io_ret_0_2 => shiftrows4_io_ret_0_2,
      io_ret_0_3 => shiftrows4_io_ret_0_3,
      io_ret_1_0 => shiftrows4_io_ret_1_0,
      io_ret_1_1 => shiftrows4_io_ret_1_1,
      io_ret_1_2 => shiftrows4_io_ret_1_2,
      io_ret_1_3 => shiftrows4_io_ret_1_3,
      io_ret_2_0 => shiftrows4_io_ret_2_0,
      io_ret_2_1 => shiftrows4_io_ret_2_1,
      io_ret_2_2 => shiftrows4_io_ret_2_2,
      io_ret_2_3 => shiftrows4_io_ret_2_3,
      io_ret_3_0 => shiftrows4_io_ret_3_0,
      io_ret_3_1 => shiftrows4_io_ret_3_1,
      io_ret_3_2 => shiftrows4_io_ret_3_2,
      io_ret_3_3 => shiftrows4_io_ret_3_3 
    );
  mixcolumns4 : entity work.MixColumns
    port map ( 
      io_state_0_0 => shiftrows4_io_ret_0_0,
      io_state_0_1 => shiftrows4_io_ret_0_1,
      io_state_0_2 => shiftrows4_io_ret_0_2,
      io_state_0_3 => shiftrows4_io_ret_0_3,
      io_state_1_0 => shiftrows4_io_ret_1_0,
      io_state_1_1 => shiftrows4_io_ret_1_1,
      io_state_1_2 => shiftrows4_io_ret_1_2,
      io_state_1_3 => shiftrows4_io_ret_1_3,
      io_state_2_0 => shiftrows4_io_ret_2_0,
      io_state_2_1 => shiftrows4_io_ret_2_1,
      io_state_2_2 => shiftrows4_io_ret_2_2,
      io_state_2_3 => shiftrows4_io_ret_2_3,
      io_state_3_0 => shiftrows4_io_ret_3_0,
      io_state_3_1 => shiftrows4_io_ret_3_1,
      io_state_3_2 => shiftrows4_io_ret_3_2,
      io_state_3_3 => shiftrows4_io_ret_3_3,
      io_ret_0_0 => mixcolumns4_io_ret_0_0,
      io_ret_0_1 => mixcolumns4_io_ret_0_1,
      io_ret_0_2 => mixcolumns4_io_ret_0_2,
      io_ret_0_3 => mixcolumns4_io_ret_0_3,
      io_ret_1_0 => mixcolumns4_io_ret_1_0,
      io_ret_1_1 => mixcolumns4_io_ret_1_1,
      io_ret_1_2 => mixcolumns4_io_ret_1_2,
      io_ret_1_3 => mixcolumns4_io_ret_1_3,
      io_ret_2_0 => mixcolumns4_io_ret_2_0,
      io_ret_2_1 => mixcolumns4_io_ret_2_1,
      io_ret_2_2 => mixcolumns4_io_ret_2_2,
      io_ret_2_3 => mixcolumns4_io_ret_2_3,
      io_ret_3_0 => mixcolumns4_io_ret_3_0,
      io_ret_3_1 => mixcolumns4_io_ret_3_1,
      io_ret_3_2 => mixcolumns4_io_ret_3_2,
      io_ret_3_3 => mixcolumns4_io_ret_3_3 
    );
  addroundkey4 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keyschedule3_io_ret_0_0,
      io_rk_0_1 => keyschedule3_io_ret_0_1,
      io_rk_0_2 => keyschedule3_io_ret_0_2,
      io_rk_0_3 => keyschedule3_io_ret_0_3,
      io_rk_1_0 => keyschedule3_io_ret_1_0,
      io_rk_1_1 => keyschedule3_io_ret_1_1,
      io_rk_1_2 => keyschedule3_io_ret_1_2,
      io_rk_1_3 => keyschedule3_io_ret_1_3,
      io_rk_2_0 => keyschedule3_io_ret_2_0,
      io_rk_2_1 => keyschedule3_io_ret_2_1,
      io_rk_2_2 => keyschedule3_io_ret_2_2,
      io_rk_2_3 => keyschedule3_io_ret_2_3,
      io_rk_3_0 => keyschedule3_io_ret_3_0,
      io_rk_3_1 => keyschedule3_io_ret_3_1,
      io_rk_3_2 => keyschedule3_io_ret_3_2,
      io_rk_3_3 => keyschedule3_io_ret_3_3,
      io_s_0_0 => mixcolumns4_io_ret_0_0,
      io_s_0_1 => mixcolumns4_io_ret_0_1,
      io_s_0_2 => mixcolumns4_io_ret_0_2,
      io_s_0_3 => mixcolumns4_io_ret_0_3,
      io_s_1_0 => mixcolumns4_io_ret_1_0,
      io_s_1_1 => mixcolumns4_io_ret_1_1,
      io_s_1_2 => mixcolumns4_io_ret_1_2,
      io_s_1_3 => mixcolumns4_io_ret_1_3,
      io_s_2_0 => mixcolumns4_io_ret_2_0,
      io_s_2_1 => mixcolumns4_io_ret_2_1,
      io_s_2_2 => mixcolumns4_io_ret_2_2,
      io_s_2_3 => mixcolumns4_io_ret_2_3,
      io_s_3_0 => mixcolumns4_io_ret_3_0,
      io_s_3_1 => mixcolumns4_io_ret_3_1,
      io_s_3_2 => mixcolumns4_io_ret_3_2,
      io_s_3_3 => mixcolumns4_io_ret_3_3,
      io_ret_0_0 => addroundkey4_io_ret_0_0,
      io_ret_0_1 => addroundkey4_io_ret_0_1,
      io_ret_0_2 => addroundkey4_io_ret_0_2,
      io_ret_0_3 => addroundkey4_io_ret_0_3,
      io_ret_1_0 => addroundkey4_io_ret_1_0,
      io_ret_1_1 => addroundkey4_io_ret_1_1,
      io_ret_1_2 => addroundkey4_io_ret_1_2,
      io_ret_1_3 => addroundkey4_io_ret_1_3,
      io_ret_2_0 => addroundkey4_io_ret_2_0,
      io_ret_2_1 => addroundkey4_io_ret_2_1,
      io_ret_2_2 => addroundkey4_io_ret_2_2,
      io_ret_2_3 => addroundkey4_io_ret_2_3,
      io_ret_3_0 => addroundkey4_io_ret_3_0,
      io_ret_3_1 => addroundkey4_io_ret_3_1,
      io_ret_3_2 => addroundkey4_io_ret_3_2,
      io_ret_3_3 => addroundkey4_io_ret_3_3 
    );
  nextrc4 : entity work.NextRC
    port map ( 
      io_rc => nextrc3_io_ret,
      io_ret => nextrc4_io_ret 
    );
  keyschedule4 : entity work.KeySchedule
    port map ( 
      io_key_0_0 => keyschedule3_io_ret_0_0,
      io_key_0_1 => keyschedule3_io_ret_0_1,
      io_key_0_2 => keyschedule3_io_ret_0_2,
      io_key_0_3 => keyschedule3_io_ret_0_3,
      io_key_1_0 => keyschedule3_io_ret_1_0,
      io_key_1_1 => keyschedule3_io_ret_1_1,
      io_key_1_2 => keyschedule3_io_ret_1_2,
      io_key_1_3 => keyschedule3_io_ret_1_3,
      io_key_2_0 => keyschedule3_io_ret_2_0,
      io_key_2_1 => keyschedule3_io_ret_2_1,
      io_key_2_2 => keyschedule3_io_ret_2_2,
      io_key_2_3 => keyschedule3_io_ret_2_3,
      io_key_3_0 => keyschedule3_io_ret_3_0,
      io_key_3_1 => keyschedule3_io_ret_3_1,
      io_key_3_2 => keyschedule3_io_ret_3_2,
      io_key_3_3 => keyschedule3_io_ret_3_3,
      io_c => nextrc3_io_ret,
      io_ret_0_0 => keyschedule4_io_ret_0_0,
      io_ret_0_1 => keyschedule4_io_ret_0_1,
      io_ret_0_2 => keyschedule4_io_ret_0_2,
      io_ret_0_3 => keyschedule4_io_ret_0_3,
      io_ret_1_0 => keyschedule4_io_ret_1_0,
      io_ret_1_1 => keyschedule4_io_ret_1_1,
      io_ret_1_2 => keyschedule4_io_ret_1_2,
      io_ret_1_3 => keyschedule4_io_ret_1_3,
      io_ret_2_0 => keyschedule4_io_ret_2_0,
      io_ret_2_1 => keyschedule4_io_ret_2_1,
      io_ret_2_2 => keyschedule4_io_ret_2_2,
      io_ret_2_3 => keyschedule4_io_ret_2_3,
      io_ret_3_0 => keyschedule4_io_ret_3_0,
      io_ret_3_1 => keyschedule4_io_ret_3_1,
      io_ret_3_2 => keyschedule4_io_ret_3_2,
      io_ret_3_3 => keyschedule4_io_ret_3_3 
    );
  subbytes5 : entity work.SubBytes
    port map ( 
      io_state_0_0 => addroundkey4_io_ret_0_0,
      io_state_0_1 => addroundkey4_io_ret_0_1,
      io_state_0_2 => addroundkey4_io_ret_0_2,
      io_state_0_3 => addroundkey4_io_ret_0_3,
      io_state_1_0 => addroundkey4_io_ret_1_0,
      io_state_1_1 => addroundkey4_io_ret_1_1,
      io_state_1_2 => addroundkey4_io_ret_1_2,
      io_state_1_3 => addroundkey4_io_ret_1_3,
      io_state_2_0 => addroundkey4_io_ret_2_0,
      io_state_2_1 => addroundkey4_io_ret_2_1,
      io_state_2_2 => addroundkey4_io_ret_2_2,
      io_state_2_3 => addroundkey4_io_ret_2_3,
      io_state_3_0 => addroundkey4_io_ret_3_0,
      io_state_3_1 => addroundkey4_io_ret_3_1,
      io_state_3_2 => addroundkey4_io_ret_3_2,
      io_state_3_3 => addroundkey4_io_ret_3_3,
      io_ret_0_0 => subbytes5_io_ret_0_0,
      io_ret_0_1 => subbytes5_io_ret_0_1,
      io_ret_0_2 => subbytes5_io_ret_0_2,
      io_ret_0_3 => subbytes5_io_ret_0_3,
      io_ret_1_0 => subbytes5_io_ret_1_0,
      io_ret_1_1 => subbytes5_io_ret_1_1,
      io_ret_1_2 => subbytes5_io_ret_1_2,
      io_ret_1_3 => subbytes5_io_ret_1_3,
      io_ret_2_0 => subbytes5_io_ret_2_0,
      io_ret_2_1 => subbytes5_io_ret_2_1,
      io_ret_2_2 => subbytes5_io_ret_2_2,
      io_ret_2_3 => subbytes5_io_ret_2_3,
      io_ret_3_0 => subbytes5_io_ret_3_0,
      io_ret_3_1 => subbytes5_io_ret_3_1,
      io_ret_3_2 => subbytes5_io_ret_3_2,
      io_ret_3_3 => subbytes5_io_ret_3_3 
    );
  shiftrows5 : entity work.ShiftRows
    port map ( 
      io_state_0_0 => subbytes5_io_ret_0_0,
      io_state_0_1 => subbytes5_io_ret_0_1,
      io_state_0_2 => subbytes5_io_ret_0_2,
      io_state_0_3 => subbytes5_io_ret_0_3,
      io_state_1_0 => subbytes5_io_ret_1_0,
      io_state_1_1 => subbytes5_io_ret_1_1,
      io_state_1_2 => subbytes5_io_ret_1_2,
      io_state_1_3 => subbytes5_io_ret_1_3,
      io_state_2_0 => subbytes5_io_ret_2_0,
      io_state_2_1 => subbytes5_io_ret_2_1,
      io_state_2_2 => subbytes5_io_ret_2_2,
      io_state_2_3 => subbytes5_io_ret_2_3,
      io_state_3_0 => subbytes5_io_ret_3_0,
      io_state_3_1 => subbytes5_io_ret_3_1,
      io_state_3_2 => subbytes5_io_ret_3_2,
      io_state_3_3 => subbytes5_io_ret_3_3,
      io_ret_0_0 => shiftrows5_io_ret_0_0,
      io_ret_0_1 => shiftrows5_io_ret_0_1,
      io_ret_0_2 => shiftrows5_io_ret_0_2,
      io_ret_0_3 => shiftrows5_io_ret_0_3,
      io_ret_1_0 => shiftrows5_io_ret_1_0,
      io_ret_1_1 => shiftrows5_io_ret_1_1,
      io_ret_1_2 => shiftrows5_io_ret_1_2,
      io_ret_1_3 => shiftrows5_io_ret_1_3,
      io_ret_2_0 => shiftrows5_io_ret_2_0,
      io_ret_2_1 => shiftrows5_io_ret_2_1,
      io_ret_2_2 => shiftrows5_io_ret_2_2,
      io_ret_2_3 => shiftrows5_io_ret_2_3,
      io_ret_3_0 => shiftrows5_io_ret_3_0,
      io_ret_3_1 => shiftrows5_io_ret_3_1,
      io_ret_3_2 => shiftrows5_io_ret_3_2,
      io_ret_3_3 => shiftrows5_io_ret_3_3 
    );
  mixcolumns5 : entity work.MixColumns
    port map ( 
      io_state_0_0 => shiftrows5_io_ret_0_0,
      io_state_0_1 => shiftrows5_io_ret_0_1,
      io_state_0_2 => shiftrows5_io_ret_0_2,
      io_state_0_3 => shiftrows5_io_ret_0_3,
      io_state_1_0 => shiftrows5_io_ret_1_0,
      io_state_1_1 => shiftrows5_io_ret_1_1,
      io_state_1_2 => shiftrows5_io_ret_1_2,
      io_state_1_3 => shiftrows5_io_ret_1_3,
      io_state_2_0 => shiftrows5_io_ret_2_0,
      io_state_2_1 => shiftrows5_io_ret_2_1,
      io_state_2_2 => shiftrows5_io_ret_2_2,
      io_state_2_3 => shiftrows5_io_ret_2_3,
      io_state_3_0 => shiftrows5_io_ret_3_0,
      io_state_3_1 => shiftrows5_io_ret_3_1,
      io_state_3_2 => shiftrows5_io_ret_3_2,
      io_state_3_3 => shiftrows5_io_ret_3_3,
      io_ret_0_0 => mixcolumns5_io_ret_0_0,
      io_ret_0_1 => mixcolumns5_io_ret_0_1,
      io_ret_0_2 => mixcolumns5_io_ret_0_2,
      io_ret_0_3 => mixcolumns5_io_ret_0_3,
      io_ret_1_0 => mixcolumns5_io_ret_1_0,
      io_ret_1_1 => mixcolumns5_io_ret_1_1,
      io_ret_1_2 => mixcolumns5_io_ret_1_2,
      io_ret_1_3 => mixcolumns5_io_ret_1_3,
      io_ret_2_0 => mixcolumns5_io_ret_2_0,
      io_ret_2_1 => mixcolumns5_io_ret_2_1,
      io_ret_2_2 => mixcolumns5_io_ret_2_2,
      io_ret_2_3 => mixcolumns5_io_ret_2_3,
      io_ret_3_0 => mixcolumns5_io_ret_3_0,
      io_ret_3_1 => mixcolumns5_io_ret_3_1,
      io_ret_3_2 => mixcolumns5_io_ret_3_2,
      io_ret_3_3 => mixcolumns5_io_ret_3_3 
    );
  addroundkey5 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keyschedule4_io_ret_0_0,
      io_rk_0_1 => keyschedule4_io_ret_0_1,
      io_rk_0_2 => keyschedule4_io_ret_0_2,
      io_rk_0_3 => keyschedule4_io_ret_0_3,
      io_rk_1_0 => keyschedule4_io_ret_1_0,
      io_rk_1_1 => keyschedule4_io_ret_1_1,
      io_rk_1_2 => keyschedule4_io_ret_1_2,
      io_rk_1_3 => keyschedule4_io_ret_1_3,
      io_rk_2_0 => keyschedule4_io_ret_2_0,
      io_rk_2_1 => keyschedule4_io_ret_2_1,
      io_rk_2_2 => keyschedule4_io_ret_2_2,
      io_rk_2_3 => keyschedule4_io_ret_2_3,
      io_rk_3_0 => keyschedule4_io_ret_3_0,
      io_rk_3_1 => keyschedule4_io_ret_3_1,
      io_rk_3_2 => keyschedule4_io_ret_3_2,
      io_rk_3_3 => keyschedule4_io_ret_3_3,
      io_s_0_0 => mixcolumns5_io_ret_0_0,
      io_s_0_1 => mixcolumns5_io_ret_0_1,
      io_s_0_2 => mixcolumns5_io_ret_0_2,
      io_s_0_3 => mixcolumns5_io_ret_0_3,
      io_s_1_0 => mixcolumns5_io_ret_1_0,
      io_s_1_1 => mixcolumns5_io_ret_1_1,
      io_s_1_2 => mixcolumns5_io_ret_1_2,
      io_s_1_3 => mixcolumns5_io_ret_1_3,
      io_s_2_0 => mixcolumns5_io_ret_2_0,
      io_s_2_1 => mixcolumns5_io_ret_2_1,
      io_s_2_2 => mixcolumns5_io_ret_2_2,
      io_s_2_3 => mixcolumns5_io_ret_2_3,
      io_s_3_0 => mixcolumns5_io_ret_3_0,
      io_s_3_1 => mixcolumns5_io_ret_3_1,
      io_s_3_2 => mixcolumns5_io_ret_3_2,
      io_s_3_3 => mixcolumns5_io_ret_3_3,
      io_ret_0_0 => addroundkey5_io_ret_0_0,
      io_ret_0_1 => addroundkey5_io_ret_0_1,
      io_ret_0_2 => addroundkey5_io_ret_0_2,
      io_ret_0_3 => addroundkey5_io_ret_0_3,
      io_ret_1_0 => addroundkey5_io_ret_1_0,
      io_ret_1_1 => addroundkey5_io_ret_1_1,
      io_ret_1_2 => addroundkey5_io_ret_1_2,
      io_ret_1_3 => addroundkey5_io_ret_1_3,
      io_ret_2_0 => addroundkey5_io_ret_2_0,
      io_ret_2_1 => addroundkey5_io_ret_2_1,
      io_ret_2_2 => addroundkey5_io_ret_2_2,
      io_ret_2_3 => addroundkey5_io_ret_2_3,
      io_ret_3_0 => addroundkey5_io_ret_3_0,
      io_ret_3_1 => addroundkey5_io_ret_3_1,
      io_ret_3_2 => addroundkey5_io_ret_3_2,
      io_ret_3_3 => addroundkey5_io_ret_3_3 
    );
  nextrc5 : entity work.NextRC
    port map ( 
      io_rc => nextrc4_io_ret,
      io_ret => nextrc5_io_ret 
    );
  keyschedule5 : entity work.KeySchedule
    port map ( 
      io_key_0_0 => keyschedule4_io_ret_0_0,
      io_key_0_1 => keyschedule4_io_ret_0_1,
      io_key_0_2 => keyschedule4_io_ret_0_2,
      io_key_0_3 => keyschedule4_io_ret_0_3,
      io_key_1_0 => keyschedule4_io_ret_1_0,
      io_key_1_1 => keyschedule4_io_ret_1_1,
      io_key_1_2 => keyschedule4_io_ret_1_2,
      io_key_1_3 => keyschedule4_io_ret_1_3,
      io_key_2_0 => keyschedule4_io_ret_2_0,
      io_key_2_1 => keyschedule4_io_ret_2_1,
      io_key_2_2 => keyschedule4_io_ret_2_2,
      io_key_2_3 => keyschedule4_io_ret_2_3,
      io_key_3_0 => keyschedule4_io_ret_3_0,
      io_key_3_1 => keyschedule4_io_ret_3_1,
      io_key_3_2 => keyschedule4_io_ret_3_2,
      io_key_3_3 => keyschedule4_io_ret_3_3,
      io_c => nextrc4_io_ret,
      io_ret_0_0 => keyschedule5_io_ret_0_0,
      io_ret_0_1 => keyschedule5_io_ret_0_1,
      io_ret_0_2 => keyschedule5_io_ret_0_2,
      io_ret_0_3 => keyschedule5_io_ret_0_3,
      io_ret_1_0 => keyschedule5_io_ret_1_0,
      io_ret_1_1 => keyschedule5_io_ret_1_1,
      io_ret_1_2 => keyschedule5_io_ret_1_2,
      io_ret_1_3 => keyschedule5_io_ret_1_3,
      io_ret_2_0 => keyschedule5_io_ret_2_0,
      io_ret_2_1 => keyschedule5_io_ret_2_1,
      io_ret_2_2 => keyschedule5_io_ret_2_2,
      io_ret_2_3 => keyschedule5_io_ret_2_3,
      io_ret_3_0 => keyschedule5_io_ret_3_0,
      io_ret_3_1 => keyschedule5_io_ret_3_1,
      io_ret_3_2 => keyschedule5_io_ret_3_2,
      io_ret_3_3 => keyschedule5_io_ret_3_3 
    );
  subbytes6 : entity work.SubBytes
    port map ( 
      io_state_0_0 => addroundkey5_io_ret_0_0,
      io_state_0_1 => addroundkey5_io_ret_0_1,
      io_state_0_2 => addroundkey5_io_ret_0_2,
      io_state_0_3 => addroundkey5_io_ret_0_3,
      io_state_1_0 => addroundkey5_io_ret_1_0,
      io_state_1_1 => addroundkey5_io_ret_1_1,
      io_state_1_2 => addroundkey5_io_ret_1_2,
      io_state_1_3 => addroundkey5_io_ret_1_3,
      io_state_2_0 => addroundkey5_io_ret_2_0,
      io_state_2_1 => addroundkey5_io_ret_2_1,
      io_state_2_2 => addroundkey5_io_ret_2_2,
      io_state_2_3 => addroundkey5_io_ret_2_3,
      io_state_3_0 => addroundkey5_io_ret_3_0,
      io_state_3_1 => addroundkey5_io_ret_3_1,
      io_state_3_2 => addroundkey5_io_ret_3_2,
      io_state_3_3 => addroundkey5_io_ret_3_3,
      io_ret_0_0 => subbytes6_io_ret_0_0,
      io_ret_0_1 => subbytes6_io_ret_0_1,
      io_ret_0_2 => subbytes6_io_ret_0_2,
      io_ret_0_3 => subbytes6_io_ret_0_3,
      io_ret_1_0 => subbytes6_io_ret_1_0,
      io_ret_1_1 => subbytes6_io_ret_1_1,
      io_ret_1_2 => subbytes6_io_ret_1_2,
      io_ret_1_3 => subbytes6_io_ret_1_3,
      io_ret_2_0 => subbytes6_io_ret_2_0,
      io_ret_2_1 => subbytes6_io_ret_2_1,
      io_ret_2_2 => subbytes6_io_ret_2_2,
      io_ret_2_3 => subbytes6_io_ret_2_3,
      io_ret_3_0 => subbytes6_io_ret_3_0,
      io_ret_3_1 => subbytes6_io_ret_3_1,
      io_ret_3_2 => subbytes6_io_ret_3_2,
      io_ret_3_3 => subbytes6_io_ret_3_3 
    );
  shiftrows6 : entity work.ShiftRows
    port map ( 
      io_state_0_0 => subbytes6_io_ret_0_0,
      io_state_0_1 => subbytes6_io_ret_0_1,
      io_state_0_2 => subbytes6_io_ret_0_2,
      io_state_0_3 => subbytes6_io_ret_0_3,
      io_state_1_0 => subbytes6_io_ret_1_0,
      io_state_1_1 => subbytes6_io_ret_1_1,
      io_state_1_2 => subbytes6_io_ret_1_2,
      io_state_1_3 => subbytes6_io_ret_1_3,
      io_state_2_0 => subbytes6_io_ret_2_0,
      io_state_2_1 => subbytes6_io_ret_2_1,
      io_state_2_2 => subbytes6_io_ret_2_2,
      io_state_2_3 => subbytes6_io_ret_2_3,
      io_state_3_0 => subbytes6_io_ret_3_0,
      io_state_3_1 => subbytes6_io_ret_3_1,
      io_state_3_2 => subbytes6_io_ret_3_2,
      io_state_3_3 => subbytes6_io_ret_3_3,
      io_ret_0_0 => shiftrows6_io_ret_0_0,
      io_ret_0_1 => shiftrows6_io_ret_0_1,
      io_ret_0_2 => shiftrows6_io_ret_0_2,
      io_ret_0_3 => shiftrows6_io_ret_0_3,
      io_ret_1_0 => shiftrows6_io_ret_1_0,
      io_ret_1_1 => shiftrows6_io_ret_1_1,
      io_ret_1_2 => shiftrows6_io_ret_1_2,
      io_ret_1_3 => shiftrows6_io_ret_1_3,
      io_ret_2_0 => shiftrows6_io_ret_2_0,
      io_ret_2_1 => shiftrows6_io_ret_2_1,
      io_ret_2_2 => shiftrows6_io_ret_2_2,
      io_ret_2_3 => shiftrows6_io_ret_2_3,
      io_ret_3_0 => shiftrows6_io_ret_3_0,
      io_ret_3_1 => shiftrows6_io_ret_3_1,
      io_ret_3_2 => shiftrows6_io_ret_3_2,
      io_ret_3_3 => shiftrows6_io_ret_3_3 
    );
  mixcolumns6 : entity work.MixColumns
    port map ( 
      io_state_0_0 => shiftrows6_io_ret_0_0,
      io_state_0_1 => shiftrows6_io_ret_0_1,
      io_state_0_2 => shiftrows6_io_ret_0_2,
      io_state_0_3 => shiftrows6_io_ret_0_3,
      io_state_1_0 => shiftrows6_io_ret_1_0,
      io_state_1_1 => shiftrows6_io_ret_1_1,
      io_state_1_2 => shiftrows6_io_ret_1_2,
      io_state_1_3 => shiftrows6_io_ret_1_3,
      io_state_2_0 => shiftrows6_io_ret_2_0,
      io_state_2_1 => shiftrows6_io_ret_2_1,
      io_state_2_2 => shiftrows6_io_ret_2_2,
      io_state_2_3 => shiftrows6_io_ret_2_3,
      io_state_3_0 => shiftrows6_io_ret_3_0,
      io_state_3_1 => shiftrows6_io_ret_3_1,
      io_state_3_2 => shiftrows6_io_ret_3_2,
      io_state_3_3 => shiftrows6_io_ret_3_3,
      io_ret_0_0 => mixcolumns6_io_ret_0_0,
      io_ret_0_1 => mixcolumns6_io_ret_0_1,
      io_ret_0_2 => mixcolumns6_io_ret_0_2,
      io_ret_0_3 => mixcolumns6_io_ret_0_3,
      io_ret_1_0 => mixcolumns6_io_ret_1_0,
      io_ret_1_1 => mixcolumns6_io_ret_1_1,
      io_ret_1_2 => mixcolumns6_io_ret_1_2,
      io_ret_1_3 => mixcolumns6_io_ret_1_3,
      io_ret_2_0 => mixcolumns6_io_ret_2_0,
      io_ret_2_1 => mixcolumns6_io_ret_2_1,
      io_ret_2_2 => mixcolumns6_io_ret_2_2,
      io_ret_2_3 => mixcolumns6_io_ret_2_3,
      io_ret_3_0 => mixcolumns6_io_ret_3_0,
      io_ret_3_1 => mixcolumns6_io_ret_3_1,
      io_ret_3_2 => mixcolumns6_io_ret_3_2,
      io_ret_3_3 => mixcolumns6_io_ret_3_3 
    );
  addroundkey6 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keyschedule5_io_ret_0_0,
      io_rk_0_1 => keyschedule5_io_ret_0_1,
      io_rk_0_2 => keyschedule5_io_ret_0_2,
      io_rk_0_3 => keyschedule5_io_ret_0_3,
      io_rk_1_0 => keyschedule5_io_ret_1_0,
      io_rk_1_1 => keyschedule5_io_ret_1_1,
      io_rk_1_2 => keyschedule5_io_ret_1_2,
      io_rk_1_3 => keyschedule5_io_ret_1_3,
      io_rk_2_0 => keyschedule5_io_ret_2_0,
      io_rk_2_1 => keyschedule5_io_ret_2_1,
      io_rk_2_2 => keyschedule5_io_ret_2_2,
      io_rk_2_3 => keyschedule5_io_ret_2_3,
      io_rk_3_0 => keyschedule5_io_ret_3_0,
      io_rk_3_1 => keyschedule5_io_ret_3_1,
      io_rk_3_2 => keyschedule5_io_ret_3_2,
      io_rk_3_3 => keyschedule5_io_ret_3_3,
      io_s_0_0 => mixcolumns6_io_ret_0_0,
      io_s_0_1 => mixcolumns6_io_ret_0_1,
      io_s_0_2 => mixcolumns6_io_ret_0_2,
      io_s_0_3 => mixcolumns6_io_ret_0_3,
      io_s_1_0 => mixcolumns6_io_ret_1_0,
      io_s_1_1 => mixcolumns6_io_ret_1_1,
      io_s_1_2 => mixcolumns6_io_ret_1_2,
      io_s_1_3 => mixcolumns6_io_ret_1_3,
      io_s_2_0 => mixcolumns6_io_ret_2_0,
      io_s_2_1 => mixcolumns6_io_ret_2_1,
      io_s_2_2 => mixcolumns6_io_ret_2_2,
      io_s_2_3 => mixcolumns6_io_ret_2_3,
      io_s_3_0 => mixcolumns6_io_ret_3_0,
      io_s_3_1 => mixcolumns6_io_ret_3_1,
      io_s_3_2 => mixcolumns6_io_ret_3_2,
      io_s_3_3 => mixcolumns6_io_ret_3_3,
      io_ret_0_0 => addroundkey6_io_ret_0_0,
      io_ret_0_1 => addroundkey6_io_ret_0_1,
      io_ret_0_2 => addroundkey6_io_ret_0_2,
      io_ret_0_3 => addroundkey6_io_ret_0_3,
      io_ret_1_0 => addroundkey6_io_ret_1_0,
      io_ret_1_1 => addroundkey6_io_ret_1_1,
      io_ret_1_2 => addroundkey6_io_ret_1_2,
      io_ret_1_3 => addroundkey6_io_ret_1_3,
      io_ret_2_0 => addroundkey6_io_ret_2_0,
      io_ret_2_1 => addroundkey6_io_ret_2_1,
      io_ret_2_2 => addroundkey6_io_ret_2_2,
      io_ret_2_3 => addroundkey6_io_ret_2_3,
      io_ret_3_0 => addroundkey6_io_ret_3_0,
      io_ret_3_1 => addroundkey6_io_ret_3_1,
      io_ret_3_2 => addroundkey6_io_ret_3_2,
      io_ret_3_3 => addroundkey6_io_ret_3_3 
    );
  nextrc6 : entity work.NextRC
    port map ( 
      io_rc => nextrc5_io_ret,
      io_ret => nextrc6_io_ret 
    );
  keyschedule6 : entity work.KeySchedule
    port map ( 
      io_key_0_0 => keyschedule5_io_ret_0_0,
      io_key_0_1 => keyschedule5_io_ret_0_1,
      io_key_0_2 => keyschedule5_io_ret_0_2,
      io_key_0_3 => keyschedule5_io_ret_0_3,
      io_key_1_0 => keyschedule5_io_ret_1_0,
      io_key_1_1 => keyschedule5_io_ret_1_1,
      io_key_1_2 => keyschedule5_io_ret_1_2,
      io_key_1_3 => keyschedule5_io_ret_1_3,
      io_key_2_0 => keyschedule5_io_ret_2_0,
      io_key_2_1 => keyschedule5_io_ret_2_1,
      io_key_2_2 => keyschedule5_io_ret_2_2,
      io_key_2_3 => keyschedule5_io_ret_2_3,
      io_key_3_0 => keyschedule5_io_ret_3_0,
      io_key_3_1 => keyschedule5_io_ret_3_1,
      io_key_3_2 => keyschedule5_io_ret_3_2,
      io_key_3_3 => keyschedule5_io_ret_3_3,
      io_c => nextrc5_io_ret,
      io_ret_0_0 => keyschedule6_io_ret_0_0,
      io_ret_0_1 => keyschedule6_io_ret_0_1,
      io_ret_0_2 => keyschedule6_io_ret_0_2,
      io_ret_0_3 => keyschedule6_io_ret_0_3,
      io_ret_1_0 => keyschedule6_io_ret_1_0,
      io_ret_1_1 => keyschedule6_io_ret_1_1,
      io_ret_1_2 => keyschedule6_io_ret_1_2,
      io_ret_1_3 => keyschedule6_io_ret_1_3,
      io_ret_2_0 => keyschedule6_io_ret_2_0,
      io_ret_2_1 => keyschedule6_io_ret_2_1,
      io_ret_2_2 => keyschedule6_io_ret_2_2,
      io_ret_2_3 => keyschedule6_io_ret_2_3,
      io_ret_3_0 => keyschedule6_io_ret_3_0,
      io_ret_3_1 => keyschedule6_io_ret_3_1,
      io_ret_3_2 => keyschedule6_io_ret_3_2,
      io_ret_3_3 => keyschedule6_io_ret_3_3 
    );
  subbytes7 : entity work.SubBytes
    port map ( 
      io_state_0_0 => addroundkey6_io_ret_0_0,
      io_state_0_1 => addroundkey6_io_ret_0_1,
      io_state_0_2 => addroundkey6_io_ret_0_2,
      io_state_0_3 => addroundkey6_io_ret_0_3,
      io_state_1_0 => addroundkey6_io_ret_1_0,
      io_state_1_1 => addroundkey6_io_ret_1_1,
      io_state_1_2 => addroundkey6_io_ret_1_2,
      io_state_1_3 => addroundkey6_io_ret_1_3,
      io_state_2_0 => addroundkey6_io_ret_2_0,
      io_state_2_1 => addroundkey6_io_ret_2_1,
      io_state_2_2 => addroundkey6_io_ret_2_2,
      io_state_2_3 => addroundkey6_io_ret_2_3,
      io_state_3_0 => addroundkey6_io_ret_3_0,
      io_state_3_1 => addroundkey6_io_ret_3_1,
      io_state_3_2 => addroundkey6_io_ret_3_2,
      io_state_3_3 => addroundkey6_io_ret_3_3,
      io_ret_0_0 => subbytes7_io_ret_0_0,
      io_ret_0_1 => subbytes7_io_ret_0_1,
      io_ret_0_2 => subbytes7_io_ret_0_2,
      io_ret_0_3 => subbytes7_io_ret_0_3,
      io_ret_1_0 => subbytes7_io_ret_1_0,
      io_ret_1_1 => subbytes7_io_ret_1_1,
      io_ret_1_2 => subbytes7_io_ret_1_2,
      io_ret_1_3 => subbytes7_io_ret_1_3,
      io_ret_2_0 => subbytes7_io_ret_2_0,
      io_ret_2_1 => subbytes7_io_ret_2_1,
      io_ret_2_2 => subbytes7_io_ret_2_2,
      io_ret_2_3 => subbytes7_io_ret_2_3,
      io_ret_3_0 => subbytes7_io_ret_3_0,
      io_ret_3_1 => subbytes7_io_ret_3_1,
      io_ret_3_2 => subbytes7_io_ret_3_2,
      io_ret_3_3 => subbytes7_io_ret_3_3 
    );
  shiftrows7 : entity work.ShiftRows
    port map ( 
      io_state_0_0 => subbytes7_io_ret_0_0,
      io_state_0_1 => subbytes7_io_ret_0_1,
      io_state_0_2 => subbytes7_io_ret_0_2,
      io_state_0_3 => subbytes7_io_ret_0_3,
      io_state_1_0 => subbytes7_io_ret_1_0,
      io_state_1_1 => subbytes7_io_ret_1_1,
      io_state_1_2 => subbytes7_io_ret_1_2,
      io_state_1_3 => subbytes7_io_ret_1_3,
      io_state_2_0 => subbytes7_io_ret_2_0,
      io_state_2_1 => subbytes7_io_ret_2_1,
      io_state_2_2 => subbytes7_io_ret_2_2,
      io_state_2_3 => subbytes7_io_ret_2_3,
      io_state_3_0 => subbytes7_io_ret_3_0,
      io_state_3_1 => subbytes7_io_ret_3_1,
      io_state_3_2 => subbytes7_io_ret_3_2,
      io_state_3_3 => subbytes7_io_ret_3_3,
      io_ret_0_0 => shiftrows7_io_ret_0_0,
      io_ret_0_1 => shiftrows7_io_ret_0_1,
      io_ret_0_2 => shiftrows7_io_ret_0_2,
      io_ret_0_3 => shiftrows7_io_ret_0_3,
      io_ret_1_0 => shiftrows7_io_ret_1_0,
      io_ret_1_1 => shiftrows7_io_ret_1_1,
      io_ret_1_2 => shiftrows7_io_ret_1_2,
      io_ret_1_3 => shiftrows7_io_ret_1_3,
      io_ret_2_0 => shiftrows7_io_ret_2_0,
      io_ret_2_1 => shiftrows7_io_ret_2_1,
      io_ret_2_2 => shiftrows7_io_ret_2_2,
      io_ret_2_3 => shiftrows7_io_ret_2_3,
      io_ret_3_0 => shiftrows7_io_ret_3_0,
      io_ret_3_1 => shiftrows7_io_ret_3_1,
      io_ret_3_2 => shiftrows7_io_ret_3_2,
      io_ret_3_3 => shiftrows7_io_ret_3_3 
    );
  mixcolumns7 : entity work.MixColumns
    port map ( 
      io_state_0_0 => shiftrows7_io_ret_0_0,
      io_state_0_1 => shiftrows7_io_ret_0_1,
      io_state_0_2 => shiftrows7_io_ret_0_2,
      io_state_0_3 => shiftrows7_io_ret_0_3,
      io_state_1_0 => shiftrows7_io_ret_1_0,
      io_state_1_1 => shiftrows7_io_ret_1_1,
      io_state_1_2 => shiftrows7_io_ret_1_2,
      io_state_1_3 => shiftrows7_io_ret_1_3,
      io_state_2_0 => shiftrows7_io_ret_2_0,
      io_state_2_1 => shiftrows7_io_ret_2_1,
      io_state_2_2 => shiftrows7_io_ret_2_2,
      io_state_2_3 => shiftrows7_io_ret_2_3,
      io_state_3_0 => shiftrows7_io_ret_3_0,
      io_state_3_1 => shiftrows7_io_ret_3_1,
      io_state_3_2 => shiftrows7_io_ret_3_2,
      io_state_3_3 => shiftrows7_io_ret_3_3,
      io_ret_0_0 => mixcolumns7_io_ret_0_0,
      io_ret_0_1 => mixcolumns7_io_ret_0_1,
      io_ret_0_2 => mixcolumns7_io_ret_0_2,
      io_ret_0_3 => mixcolumns7_io_ret_0_3,
      io_ret_1_0 => mixcolumns7_io_ret_1_0,
      io_ret_1_1 => mixcolumns7_io_ret_1_1,
      io_ret_1_2 => mixcolumns7_io_ret_1_2,
      io_ret_1_3 => mixcolumns7_io_ret_1_3,
      io_ret_2_0 => mixcolumns7_io_ret_2_0,
      io_ret_2_1 => mixcolumns7_io_ret_2_1,
      io_ret_2_2 => mixcolumns7_io_ret_2_2,
      io_ret_2_3 => mixcolumns7_io_ret_2_3,
      io_ret_3_0 => mixcolumns7_io_ret_3_0,
      io_ret_3_1 => mixcolumns7_io_ret_3_1,
      io_ret_3_2 => mixcolumns7_io_ret_3_2,
      io_ret_3_3 => mixcolumns7_io_ret_3_3 
    );
  addroundkey7 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keyschedule6_io_ret_0_0,
      io_rk_0_1 => keyschedule6_io_ret_0_1,
      io_rk_0_2 => keyschedule6_io_ret_0_2,
      io_rk_0_3 => keyschedule6_io_ret_0_3,
      io_rk_1_0 => keyschedule6_io_ret_1_0,
      io_rk_1_1 => keyschedule6_io_ret_1_1,
      io_rk_1_2 => keyschedule6_io_ret_1_2,
      io_rk_1_3 => keyschedule6_io_ret_1_3,
      io_rk_2_0 => keyschedule6_io_ret_2_0,
      io_rk_2_1 => keyschedule6_io_ret_2_1,
      io_rk_2_2 => keyschedule6_io_ret_2_2,
      io_rk_2_3 => keyschedule6_io_ret_2_3,
      io_rk_3_0 => keyschedule6_io_ret_3_0,
      io_rk_3_1 => keyschedule6_io_ret_3_1,
      io_rk_3_2 => keyschedule6_io_ret_3_2,
      io_rk_3_3 => keyschedule6_io_ret_3_3,
      io_s_0_0 => mixcolumns7_io_ret_0_0,
      io_s_0_1 => mixcolumns7_io_ret_0_1,
      io_s_0_2 => mixcolumns7_io_ret_0_2,
      io_s_0_3 => mixcolumns7_io_ret_0_3,
      io_s_1_0 => mixcolumns7_io_ret_1_0,
      io_s_1_1 => mixcolumns7_io_ret_1_1,
      io_s_1_2 => mixcolumns7_io_ret_1_2,
      io_s_1_3 => mixcolumns7_io_ret_1_3,
      io_s_2_0 => mixcolumns7_io_ret_2_0,
      io_s_2_1 => mixcolumns7_io_ret_2_1,
      io_s_2_2 => mixcolumns7_io_ret_2_2,
      io_s_2_3 => mixcolumns7_io_ret_2_3,
      io_s_3_0 => mixcolumns7_io_ret_3_0,
      io_s_3_1 => mixcolumns7_io_ret_3_1,
      io_s_3_2 => mixcolumns7_io_ret_3_2,
      io_s_3_3 => mixcolumns7_io_ret_3_3,
      io_ret_0_0 => addroundkey7_io_ret_0_0,
      io_ret_0_1 => addroundkey7_io_ret_0_1,
      io_ret_0_2 => addroundkey7_io_ret_0_2,
      io_ret_0_3 => addroundkey7_io_ret_0_3,
      io_ret_1_0 => addroundkey7_io_ret_1_0,
      io_ret_1_1 => addroundkey7_io_ret_1_1,
      io_ret_1_2 => addroundkey7_io_ret_1_2,
      io_ret_1_3 => addroundkey7_io_ret_1_3,
      io_ret_2_0 => addroundkey7_io_ret_2_0,
      io_ret_2_1 => addroundkey7_io_ret_2_1,
      io_ret_2_2 => addroundkey7_io_ret_2_2,
      io_ret_2_3 => addroundkey7_io_ret_2_3,
      io_ret_3_0 => addroundkey7_io_ret_3_0,
      io_ret_3_1 => addroundkey7_io_ret_3_1,
      io_ret_3_2 => addroundkey7_io_ret_3_2,
      io_ret_3_3 => addroundkey7_io_ret_3_3 
    );
  nextrc7 : entity work.NextRC
    port map ( 
      io_rc => nextrc6_io_ret,
      io_ret => nextrc7_io_ret 
    );
  keyschedule7 : entity work.KeySchedule
    port map ( 
      io_key_0_0 => keyschedule6_io_ret_0_0,
      io_key_0_1 => keyschedule6_io_ret_0_1,
      io_key_0_2 => keyschedule6_io_ret_0_2,
      io_key_0_3 => keyschedule6_io_ret_0_3,
      io_key_1_0 => keyschedule6_io_ret_1_0,
      io_key_1_1 => keyschedule6_io_ret_1_1,
      io_key_1_2 => keyschedule6_io_ret_1_2,
      io_key_1_3 => keyschedule6_io_ret_1_3,
      io_key_2_0 => keyschedule6_io_ret_2_0,
      io_key_2_1 => keyschedule6_io_ret_2_1,
      io_key_2_2 => keyschedule6_io_ret_2_2,
      io_key_2_3 => keyschedule6_io_ret_2_3,
      io_key_3_0 => keyschedule6_io_ret_3_0,
      io_key_3_1 => keyschedule6_io_ret_3_1,
      io_key_3_2 => keyschedule6_io_ret_3_2,
      io_key_3_3 => keyschedule6_io_ret_3_3,
      io_c => nextrc6_io_ret,
      io_ret_0_0 => keyschedule7_io_ret_0_0,
      io_ret_0_1 => keyschedule7_io_ret_0_1,
      io_ret_0_2 => keyschedule7_io_ret_0_2,
      io_ret_0_3 => keyschedule7_io_ret_0_3,
      io_ret_1_0 => keyschedule7_io_ret_1_0,
      io_ret_1_1 => keyschedule7_io_ret_1_1,
      io_ret_1_2 => keyschedule7_io_ret_1_2,
      io_ret_1_3 => keyschedule7_io_ret_1_3,
      io_ret_2_0 => keyschedule7_io_ret_2_0,
      io_ret_2_1 => keyschedule7_io_ret_2_1,
      io_ret_2_2 => keyschedule7_io_ret_2_2,
      io_ret_2_3 => keyschedule7_io_ret_2_3,
      io_ret_3_0 => keyschedule7_io_ret_3_0,
      io_ret_3_1 => keyschedule7_io_ret_3_1,
      io_ret_3_2 => keyschedule7_io_ret_3_2,
      io_ret_3_3 => keyschedule7_io_ret_3_3 
    );
  subbytes8 : entity work.SubBytes
    port map ( 
      io_state_0_0 => addroundkey7_io_ret_0_0,
      io_state_0_1 => addroundkey7_io_ret_0_1,
      io_state_0_2 => addroundkey7_io_ret_0_2,
      io_state_0_3 => addroundkey7_io_ret_0_3,
      io_state_1_0 => addroundkey7_io_ret_1_0,
      io_state_1_1 => addroundkey7_io_ret_1_1,
      io_state_1_2 => addroundkey7_io_ret_1_2,
      io_state_1_3 => addroundkey7_io_ret_1_3,
      io_state_2_0 => addroundkey7_io_ret_2_0,
      io_state_2_1 => addroundkey7_io_ret_2_1,
      io_state_2_2 => addroundkey7_io_ret_2_2,
      io_state_2_3 => addroundkey7_io_ret_2_3,
      io_state_3_0 => addroundkey7_io_ret_3_0,
      io_state_3_1 => addroundkey7_io_ret_3_1,
      io_state_3_2 => addroundkey7_io_ret_3_2,
      io_state_3_3 => addroundkey7_io_ret_3_3,
      io_ret_0_0 => subbytes8_io_ret_0_0,
      io_ret_0_1 => subbytes8_io_ret_0_1,
      io_ret_0_2 => subbytes8_io_ret_0_2,
      io_ret_0_3 => subbytes8_io_ret_0_3,
      io_ret_1_0 => subbytes8_io_ret_1_0,
      io_ret_1_1 => subbytes8_io_ret_1_1,
      io_ret_1_2 => subbytes8_io_ret_1_2,
      io_ret_1_3 => subbytes8_io_ret_1_3,
      io_ret_2_0 => subbytes8_io_ret_2_0,
      io_ret_2_1 => subbytes8_io_ret_2_1,
      io_ret_2_2 => subbytes8_io_ret_2_2,
      io_ret_2_3 => subbytes8_io_ret_2_3,
      io_ret_3_0 => subbytes8_io_ret_3_0,
      io_ret_3_1 => subbytes8_io_ret_3_1,
      io_ret_3_2 => subbytes8_io_ret_3_2,
      io_ret_3_3 => subbytes8_io_ret_3_3 
    );
  shiftrows8 : entity work.ShiftRows
    port map ( 
      io_state_0_0 => subbytes8_io_ret_0_0,
      io_state_0_1 => subbytes8_io_ret_0_1,
      io_state_0_2 => subbytes8_io_ret_0_2,
      io_state_0_3 => subbytes8_io_ret_0_3,
      io_state_1_0 => subbytes8_io_ret_1_0,
      io_state_1_1 => subbytes8_io_ret_1_1,
      io_state_1_2 => subbytes8_io_ret_1_2,
      io_state_1_3 => subbytes8_io_ret_1_3,
      io_state_2_0 => subbytes8_io_ret_2_0,
      io_state_2_1 => subbytes8_io_ret_2_1,
      io_state_2_2 => subbytes8_io_ret_2_2,
      io_state_2_3 => subbytes8_io_ret_2_3,
      io_state_3_0 => subbytes8_io_ret_3_0,
      io_state_3_1 => subbytes8_io_ret_3_1,
      io_state_3_2 => subbytes8_io_ret_3_2,
      io_state_3_3 => subbytes8_io_ret_3_3,
      io_ret_0_0 => shiftrows8_io_ret_0_0,
      io_ret_0_1 => shiftrows8_io_ret_0_1,
      io_ret_0_2 => shiftrows8_io_ret_0_2,
      io_ret_0_3 => shiftrows8_io_ret_0_3,
      io_ret_1_0 => shiftrows8_io_ret_1_0,
      io_ret_1_1 => shiftrows8_io_ret_1_1,
      io_ret_1_2 => shiftrows8_io_ret_1_2,
      io_ret_1_3 => shiftrows8_io_ret_1_3,
      io_ret_2_0 => shiftrows8_io_ret_2_0,
      io_ret_2_1 => shiftrows8_io_ret_2_1,
      io_ret_2_2 => shiftrows8_io_ret_2_2,
      io_ret_2_3 => shiftrows8_io_ret_2_3,
      io_ret_3_0 => shiftrows8_io_ret_3_0,
      io_ret_3_1 => shiftrows8_io_ret_3_1,
      io_ret_3_2 => shiftrows8_io_ret_3_2,
      io_ret_3_3 => shiftrows8_io_ret_3_3 
    );
  mixcolumns8 : entity work.MixColumns
    port map ( 
      io_state_0_0 => shiftrows8_io_ret_0_0,
      io_state_0_1 => shiftrows8_io_ret_0_1,
      io_state_0_2 => shiftrows8_io_ret_0_2,
      io_state_0_3 => shiftrows8_io_ret_0_3,
      io_state_1_0 => shiftrows8_io_ret_1_0,
      io_state_1_1 => shiftrows8_io_ret_1_1,
      io_state_1_2 => shiftrows8_io_ret_1_2,
      io_state_1_3 => shiftrows8_io_ret_1_3,
      io_state_2_0 => shiftrows8_io_ret_2_0,
      io_state_2_1 => shiftrows8_io_ret_2_1,
      io_state_2_2 => shiftrows8_io_ret_2_2,
      io_state_2_3 => shiftrows8_io_ret_2_3,
      io_state_3_0 => shiftrows8_io_ret_3_0,
      io_state_3_1 => shiftrows8_io_ret_3_1,
      io_state_3_2 => shiftrows8_io_ret_3_2,
      io_state_3_3 => shiftrows8_io_ret_3_3,
      io_ret_0_0 => mixcolumns8_io_ret_0_0,
      io_ret_0_1 => mixcolumns8_io_ret_0_1,
      io_ret_0_2 => mixcolumns8_io_ret_0_2,
      io_ret_0_3 => mixcolumns8_io_ret_0_3,
      io_ret_1_0 => mixcolumns8_io_ret_1_0,
      io_ret_1_1 => mixcolumns8_io_ret_1_1,
      io_ret_1_2 => mixcolumns8_io_ret_1_2,
      io_ret_1_3 => mixcolumns8_io_ret_1_3,
      io_ret_2_0 => mixcolumns8_io_ret_2_0,
      io_ret_2_1 => mixcolumns8_io_ret_2_1,
      io_ret_2_2 => mixcolumns8_io_ret_2_2,
      io_ret_2_3 => mixcolumns8_io_ret_2_3,
      io_ret_3_0 => mixcolumns8_io_ret_3_0,
      io_ret_3_1 => mixcolumns8_io_ret_3_1,
      io_ret_3_2 => mixcolumns8_io_ret_3_2,
      io_ret_3_3 => mixcolumns8_io_ret_3_3 
    );
  addroundkey8 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keyschedule7_io_ret_0_0,
      io_rk_0_1 => keyschedule7_io_ret_0_1,
      io_rk_0_2 => keyschedule7_io_ret_0_2,
      io_rk_0_3 => keyschedule7_io_ret_0_3,
      io_rk_1_0 => keyschedule7_io_ret_1_0,
      io_rk_1_1 => keyschedule7_io_ret_1_1,
      io_rk_1_2 => keyschedule7_io_ret_1_2,
      io_rk_1_3 => keyschedule7_io_ret_1_3,
      io_rk_2_0 => keyschedule7_io_ret_2_0,
      io_rk_2_1 => keyschedule7_io_ret_2_1,
      io_rk_2_2 => keyschedule7_io_ret_2_2,
      io_rk_2_3 => keyschedule7_io_ret_2_3,
      io_rk_3_0 => keyschedule7_io_ret_3_0,
      io_rk_3_1 => keyschedule7_io_ret_3_1,
      io_rk_3_2 => keyschedule7_io_ret_3_2,
      io_rk_3_3 => keyschedule7_io_ret_3_3,
      io_s_0_0 => mixcolumns8_io_ret_0_0,
      io_s_0_1 => mixcolumns8_io_ret_0_1,
      io_s_0_2 => mixcolumns8_io_ret_0_2,
      io_s_0_3 => mixcolumns8_io_ret_0_3,
      io_s_1_0 => mixcolumns8_io_ret_1_0,
      io_s_1_1 => mixcolumns8_io_ret_1_1,
      io_s_1_2 => mixcolumns8_io_ret_1_2,
      io_s_1_3 => mixcolumns8_io_ret_1_3,
      io_s_2_0 => mixcolumns8_io_ret_2_0,
      io_s_2_1 => mixcolumns8_io_ret_2_1,
      io_s_2_2 => mixcolumns8_io_ret_2_2,
      io_s_2_3 => mixcolumns8_io_ret_2_3,
      io_s_3_0 => mixcolumns8_io_ret_3_0,
      io_s_3_1 => mixcolumns8_io_ret_3_1,
      io_s_3_2 => mixcolumns8_io_ret_3_2,
      io_s_3_3 => mixcolumns8_io_ret_3_3,
      io_ret_0_0 => addroundkey8_io_ret_0_0,
      io_ret_0_1 => addroundkey8_io_ret_0_1,
      io_ret_0_2 => addroundkey8_io_ret_0_2,
      io_ret_0_3 => addroundkey8_io_ret_0_3,
      io_ret_1_0 => addroundkey8_io_ret_1_0,
      io_ret_1_1 => addroundkey8_io_ret_1_1,
      io_ret_1_2 => addroundkey8_io_ret_1_2,
      io_ret_1_3 => addroundkey8_io_ret_1_3,
      io_ret_2_0 => addroundkey8_io_ret_2_0,
      io_ret_2_1 => addroundkey8_io_ret_2_1,
      io_ret_2_2 => addroundkey8_io_ret_2_2,
      io_ret_2_3 => addroundkey8_io_ret_2_3,
      io_ret_3_0 => addroundkey8_io_ret_3_0,
      io_ret_3_1 => addroundkey8_io_ret_3_1,
      io_ret_3_2 => addroundkey8_io_ret_3_2,
      io_ret_3_3 => addroundkey8_io_ret_3_3 
    );
  nextrc8 : entity work.NextRC
    port map ( 
      io_rc => nextrc7_io_ret,
      io_ret => nextrc8_io_ret 
    );
  keyschedule8 : entity work.KeySchedule
    port map ( 
      io_key_0_0 => keyschedule7_io_ret_0_0,
      io_key_0_1 => keyschedule7_io_ret_0_1,
      io_key_0_2 => keyschedule7_io_ret_0_2,
      io_key_0_3 => keyschedule7_io_ret_0_3,
      io_key_1_0 => keyschedule7_io_ret_1_0,
      io_key_1_1 => keyschedule7_io_ret_1_1,
      io_key_1_2 => keyschedule7_io_ret_1_2,
      io_key_1_3 => keyschedule7_io_ret_1_3,
      io_key_2_0 => keyschedule7_io_ret_2_0,
      io_key_2_1 => keyschedule7_io_ret_2_1,
      io_key_2_2 => keyschedule7_io_ret_2_2,
      io_key_2_3 => keyschedule7_io_ret_2_3,
      io_key_3_0 => keyschedule7_io_ret_3_0,
      io_key_3_1 => keyschedule7_io_ret_3_1,
      io_key_3_2 => keyschedule7_io_ret_3_2,
      io_key_3_3 => keyschedule7_io_ret_3_3,
      io_c => nextrc7_io_ret,
      io_ret_0_0 => keyschedule8_io_ret_0_0,
      io_ret_0_1 => keyschedule8_io_ret_0_1,
      io_ret_0_2 => keyschedule8_io_ret_0_2,
      io_ret_0_3 => keyschedule8_io_ret_0_3,
      io_ret_1_0 => keyschedule8_io_ret_1_0,
      io_ret_1_1 => keyschedule8_io_ret_1_1,
      io_ret_1_2 => keyschedule8_io_ret_1_2,
      io_ret_1_3 => keyschedule8_io_ret_1_3,
      io_ret_2_0 => keyschedule8_io_ret_2_0,
      io_ret_2_1 => keyschedule8_io_ret_2_1,
      io_ret_2_2 => keyschedule8_io_ret_2_2,
      io_ret_2_3 => keyschedule8_io_ret_2_3,
      io_ret_3_0 => keyschedule8_io_ret_3_0,
      io_ret_3_1 => keyschedule8_io_ret_3_1,
      io_ret_3_2 => keyschedule8_io_ret_3_2,
      io_ret_3_3 => keyschedule8_io_ret_3_3 
    );
  subbytes9 : entity work.SubBytes
    port map ( 
      io_state_0_0 => addroundkey8_io_ret_0_0,
      io_state_0_1 => addroundkey8_io_ret_0_1,
      io_state_0_2 => addroundkey8_io_ret_0_2,
      io_state_0_3 => addroundkey8_io_ret_0_3,
      io_state_1_0 => addroundkey8_io_ret_1_0,
      io_state_1_1 => addroundkey8_io_ret_1_1,
      io_state_1_2 => addroundkey8_io_ret_1_2,
      io_state_1_3 => addroundkey8_io_ret_1_3,
      io_state_2_0 => addroundkey8_io_ret_2_0,
      io_state_2_1 => addroundkey8_io_ret_2_1,
      io_state_2_2 => addroundkey8_io_ret_2_2,
      io_state_2_3 => addroundkey8_io_ret_2_3,
      io_state_3_0 => addroundkey8_io_ret_3_0,
      io_state_3_1 => addroundkey8_io_ret_3_1,
      io_state_3_2 => addroundkey8_io_ret_3_2,
      io_state_3_3 => addroundkey8_io_ret_3_3,
      io_ret_0_0 => subbytes9_io_ret_0_0,
      io_ret_0_1 => subbytes9_io_ret_0_1,
      io_ret_0_2 => subbytes9_io_ret_0_2,
      io_ret_0_3 => subbytes9_io_ret_0_3,
      io_ret_1_0 => subbytes9_io_ret_1_0,
      io_ret_1_1 => subbytes9_io_ret_1_1,
      io_ret_1_2 => subbytes9_io_ret_1_2,
      io_ret_1_3 => subbytes9_io_ret_1_3,
      io_ret_2_0 => subbytes9_io_ret_2_0,
      io_ret_2_1 => subbytes9_io_ret_2_1,
      io_ret_2_2 => subbytes9_io_ret_2_2,
      io_ret_2_3 => subbytes9_io_ret_2_3,
      io_ret_3_0 => subbytes9_io_ret_3_0,
      io_ret_3_1 => subbytes9_io_ret_3_1,
      io_ret_3_2 => subbytes9_io_ret_3_2,
      io_ret_3_3 => subbytes9_io_ret_3_3 
    );
  shiftrows9 : entity work.ShiftRows
    port map ( 
      io_state_0_0 => subbytes9_io_ret_0_0,
      io_state_0_1 => subbytes9_io_ret_0_1,
      io_state_0_2 => subbytes9_io_ret_0_2,
      io_state_0_3 => subbytes9_io_ret_0_3,
      io_state_1_0 => subbytes9_io_ret_1_0,
      io_state_1_1 => subbytes9_io_ret_1_1,
      io_state_1_2 => subbytes9_io_ret_1_2,
      io_state_1_3 => subbytes9_io_ret_1_3,
      io_state_2_0 => subbytes9_io_ret_2_0,
      io_state_2_1 => subbytes9_io_ret_2_1,
      io_state_2_2 => subbytes9_io_ret_2_2,
      io_state_2_3 => subbytes9_io_ret_2_3,
      io_state_3_0 => subbytes9_io_ret_3_0,
      io_state_3_1 => subbytes9_io_ret_3_1,
      io_state_3_2 => subbytes9_io_ret_3_2,
      io_state_3_3 => subbytes9_io_ret_3_3,
      io_ret_0_0 => shiftrows9_io_ret_0_0,
      io_ret_0_1 => shiftrows9_io_ret_0_1,
      io_ret_0_2 => shiftrows9_io_ret_0_2,
      io_ret_0_3 => shiftrows9_io_ret_0_3,
      io_ret_1_0 => shiftrows9_io_ret_1_0,
      io_ret_1_1 => shiftrows9_io_ret_1_1,
      io_ret_1_2 => shiftrows9_io_ret_1_2,
      io_ret_1_3 => shiftrows9_io_ret_1_3,
      io_ret_2_0 => shiftrows9_io_ret_2_0,
      io_ret_2_1 => shiftrows9_io_ret_2_1,
      io_ret_2_2 => shiftrows9_io_ret_2_2,
      io_ret_2_3 => shiftrows9_io_ret_2_3,
      io_ret_3_0 => shiftrows9_io_ret_3_0,
      io_ret_3_1 => shiftrows9_io_ret_3_1,
      io_ret_3_2 => shiftrows9_io_ret_3_2,
      io_ret_3_3 => shiftrows9_io_ret_3_3 
    );
  mixcolumns9 : entity work.MixColumns
    port map ( 
      io_state_0_0 => shiftrows9_io_ret_0_0,
      io_state_0_1 => shiftrows9_io_ret_0_1,
      io_state_0_2 => shiftrows9_io_ret_0_2,
      io_state_0_3 => shiftrows9_io_ret_0_3,
      io_state_1_0 => shiftrows9_io_ret_1_0,
      io_state_1_1 => shiftrows9_io_ret_1_1,
      io_state_1_2 => shiftrows9_io_ret_1_2,
      io_state_1_3 => shiftrows9_io_ret_1_3,
      io_state_2_0 => shiftrows9_io_ret_2_0,
      io_state_2_1 => shiftrows9_io_ret_2_1,
      io_state_2_2 => shiftrows9_io_ret_2_2,
      io_state_2_3 => shiftrows9_io_ret_2_3,
      io_state_3_0 => shiftrows9_io_ret_3_0,
      io_state_3_1 => shiftrows9_io_ret_3_1,
      io_state_3_2 => shiftrows9_io_ret_3_2,
      io_state_3_3 => shiftrows9_io_ret_3_3,
      io_ret_0_0 => mixcolumns9_io_ret_0_0,
      io_ret_0_1 => mixcolumns9_io_ret_0_1,
      io_ret_0_2 => mixcolumns9_io_ret_0_2,
      io_ret_0_3 => mixcolumns9_io_ret_0_3,
      io_ret_1_0 => mixcolumns9_io_ret_1_0,
      io_ret_1_1 => mixcolumns9_io_ret_1_1,
      io_ret_1_2 => mixcolumns9_io_ret_1_2,
      io_ret_1_3 => mixcolumns9_io_ret_1_3,
      io_ret_2_0 => mixcolumns9_io_ret_2_0,
      io_ret_2_1 => mixcolumns9_io_ret_2_1,
      io_ret_2_2 => mixcolumns9_io_ret_2_2,
      io_ret_2_3 => mixcolumns9_io_ret_2_3,
      io_ret_3_0 => mixcolumns9_io_ret_3_0,
      io_ret_3_1 => mixcolumns9_io_ret_3_1,
      io_ret_3_2 => mixcolumns9_io_ret_3_2,
      io_ret_3_3 => mixcolumns9_io_ret_3_3 
    );
  addroundkey9 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keyschedule8_io_ret_0_0,
      io_rk_0_1 => keyschedule8_io_ret_0_1,
      io_rk_0_2 => keyschedule8_io_ret_0_2,
      io_rk_0_3 => keyschedule8_io_ret_0_3,
      io_rk_1_0 => keyschedule8_io_ret_1_0,
      io_rk_1_1 => keyschedule8_io_ret_1_1,
      io_rk_1_2 => keyschedule8_io_ret_1_2,
      io_rk_1_3 => keyschedule8_io_ret_1_3,
      io_rk_2_0 => keyschedule8_io_ret_2_0,
      io_rk_2_1 => keyschedule8_io_ret_2_1,
      io_rk_2_2 => keyschedule8_io_ret_2_2,
      io_rk_2_3 => keyschedule8_io_ret_2_3,
      io_rk_3_0 => keyschedule8_io_ret_3_0,
      io_rk_3_1 => keyschedule8_io_ret_3_1,
      io_rk_3_2 => keyschedule8_io_ret_3_2,
      io_rk_3_3 => keyschedule8_io_ret_3_3,
      io_s_0_0 => mixcolumns9_io_ret_0_0,
      io_s_0_1 => mixcolumns9_io_ret_0_1,
      io_s_0_2 => mixcolumns9_io_ret_0_2,
      io_s_0_3 => mixcolumns9_io_ret_0_3,
      io_s_1_0 => mixcolumns9_io_ret_1_0,
      io_s_1_1 => mixcolumns9_io_ret_1_1,
      io_s_1_2 => mixcolumns9_io_ret_1_2,
      io_s_1_3 => mixcolumns9_io_ret_1_3,
      io_s_2_0 => mixcolumns9_io_ret_2_0,
      io_s_2_1 => mixcolumns9_io_ret_2_1,
      io_s_2_2 => mixcolumns9_io_ret_2_2,
      io_s_2_3 => mixcolumns9_io_ret_2_3,
      io_s_3_0 => mixcolumns9_io_ret_3_0,
      io_s_3_1 => mixcolumns9_io_ret_3_1,
      io_s_3_2 => mixcolumns9_io_ret_3_2,
      io_s_3_3 => mixcolumns9_io_ret_3_3,
      io_ret_0_0 => addroundkey9_io_ret_0_0,
      io_ret_0_1 => addroundkey9_io_ret_0_1,
      io_ret_0_2 => addroundkey9_io_ret_0_2,
      io_ret_0_3 => addroundkey9_io_ret_0_3,
      io_ret_1_0 => addroundkey9_io_ret_1_0,
      io_ret_1_1 => addroundkey9_io_ret_1_1,
      io_ret_1_2 => addroundkey9_io_ret_1_2,
      io_ret_1_3 => addroundkey9_io_ret_1_3,
      io_ret_2_0 => addroundkey9_io_ret_2_0,
      io_ret_2_1 => addroundkey9_io_ret_2_1,
      io_ret_2_2 => addroundkey9_io_ret_2_2,
      io_ret_2_3 => addroundkey9_io_ret_2_3,
      io_ret_3_0 => addroundkey9_io_ret_3_0,
      io_ret_3_1 => addroundkey9_io_ret_3_1,
      io_ret_3_2 => addroundkey9_io_ret_3_2,
      io_ret_3_3 => addroundkey9_io_ret_3_3 
    );
  nextrc9 : entity work.NextRC
    port map ( 
      io_rc => nextrc8_io_ret,
      io_ret => nextrc9_io_ret 
    );
  keyschedule9 : entity work.KeySchedule
    port map ( 
      io_key_0_0 => keyschedule8_io_ret_0_0,
      io_key_0_1 => keyschedule8_io_ret_0_1,
      io_key_0_2 => keyschedule8_io_ret_0_2,
      io_key_0_3 => keyschedule8_io_ret_0_3,
      io_key_1_0 => keyschedule8_io_ret_1_0,
      io_key_1_1 => keyschedule8_io_ret_1_1,
      io_key_1_2 => keyschedule8_io_ret_1_2,
      io_key_1_3 => keyschedule8_io_ret_1_3,
      io_key_2_0 => keyschedule8_io_ret_2_0,
      io_key_2_1 => keyschedule8_io_ret_2_1,
      io_key_2_2 => keyschedule8_io_ret_2_2,
      io_key_2_3 => keyschedule8_io_ret_2_3,
      io_key_3_0 => keyschedule8_io_ret_3_0,
      io_key_3_1 => keyschedule8_io_ret_3_1,
      io_key_3_2 => keyschedule8_io_ret_3_2,
      io_key_3_3 => keyschedule8_io_ret_3_3,
      io_c => nextrc8_io_ret,
      io_ret_0_0 => keyschedule9_io_ret_0_0,
      io_ret_0_1 => keyschedule9_io_ret_0_1,
      io_ret_0_2 => keyschedule9_io_ret_0_2,
      io_ret_0_3 => keyschedule9_io_ret_0_3,
      io_ret_1_0 => keyschedule9_io_ret_1_0,
      io_ret_1_1 => keyschedule9_io_ret_1_1,
      io_ret_1_2 => keyschedule9_io_ret_1_2,
      io_ret_1_3 => keyschedule9_io_ret_1_3,
      io_ret_2_0 => keyschedule9_io_ret_2_0,
      io_ret_2_1 => keyschedule9_io_ret_2_1,
      io_ret_2_2 => keyschedule9_io_ret_2_2,
      io_ret_2_3 => keyschedule9_io_ret_2_3,
      io_ret_3_0 => keyschedule9_io_ret_3_0,
      io_ret_3_1 => keyschedule9_io_ret_3_1,
      io_ret_3_2 => keyschedule9_io_ret_3_2,
      io_ret_3_3 => keyschedule9_io_ret_3_3 
    );
  subbytes10 : entity work.SubBytes
    port map ( 
      io_state_0_0 => addroundkey9_io_ret_0_0,
      io_state_0_1 => addroundkey9_io_ret_0_1,
      io_state_0_2 => addroundkey9_io_ret_0_2,
      io_state_0_3 => addroundkey9_io_ret_0_3,
      io_state_1_0 => addroundkey9_io_ret_1_0,
      io_state_1_1 => addroundkey9_io_ret_1_1,
      io_state_1_2 => addroundkey9_io_ret_1_2,
      io_state_1_3 => addroundkey9_io_ret_1_3,
      io_state_2_0 => addroundkey9_io_ret_2_0,
      io_state_2_1 => addroundkey9_io_ret_2_1,
      io_state_2_2 => addroundkey9_io_ret_2_2,
      io_state_2_3 => addroundkey9_io_ret_2_3,
      io_state_3_0 => addroundkey9_io_ret_3_0,
      io_state_3_1 => addroundkey9_io_ret_3_1,
      io_state_3_2 => addroundkey9_io_ret_3_2,
      io_state_3_3 => addroundkey9_io_ret_3_3,
      io_ret_0_0 => subbytes10_io_ret_0_0,
      io_ret_0_1 => subbytes10_io_ret_0_1,
      io_ret_0_2 => subbytes10_io_ret_0_2,
      io_ret_0_3 => subbytes10_io_ret_0_3,
      io_ret_1_0 => subbytes10_io_ret_1_0,
      io_ret_1_1 => subbytes10_io_ret_1_1,
      io_ret_1_2 => subbytes10_io_ret_1_2,
      io_ret_1_3 => subbytes10_io_ret_1_3,
      io_ret_2_0 => subbytes10_io_ret_2_0,
      io_ret_2_1 => subbytes10_io_ret_2_1,
      io_ret_2_2 => subbytes10_io_ret_2_2,
      io_ret_2_3 => subbytes10_io_ret_2_3,
      io_ret_3_0 => subbytes10_io_ret_3_0,
      io_ret_3_1 => subbytes10_io_ret_3_1,
      io_ret_3_2 => subbytes10_io_ret_3_2,
      io_ret_3_3 => subbytes10_io_ret_3_3 
    );
  shiftrows10 : entity work.ShiftRows
    port map ( 
      io_state_0_0 => subbytes10_io_ret_0_0,
      io_state_0_1 => subbytes10_io_ret_0_1,
      io_state_0_2 => subbytes10_io_ret_0_2,
      io_state_0_3 => subbytes10_io_ret_0_3,
      io_state_1_0 => subbytes10_io_ret_1_0,
      io_state_1_1 => subbytes10_io_ret_1_1,
      io_state_1_2 => subbytes10_io_ret_1_2,
      io_state_1_3 => subbytes10_io_ret_1_3,
      io_state_2_0 => subbytes10_io_ret_2_0,
      io_state_2_1 => subbytes10_io_ret_2_1,
      io_state_2_2 => subbytes10_io_ret_2_2,
      io_state_2_3 => subbytes10_io_ret_2_3,
      io_state_3_0 => subbytes10_io_ret_3_0,
      io_state_3_1 => subbytes10_io_ret_3_1,
      io_state_3_2 => subbytes10_io_ret_3_2,
      io_state_3_3 => subbytes10_io_ret_3_3,
      io_ret_0_0 => shiftrows10_io_ret_0_0,
      io_ret_0_1 => shiftrows10_io_ret_0_1,
      io_ret_0_2 => shiftrows10_io_ret_0_2,
      io_ret_0_3 => shiftrows10_io_ret_0_3,
      io_ret_1_0 => shiftrows10_io_ret_1_0,
      io_ret_1_1 => shiftrows10_io_ret_1_1,
      io_ret_1_2 => shiftrows10_io_ret_1_2,
      io_ret_1_3 => shiftrows10_io_ret_1_3,
      io_ret_2_0 => shiftrows10_io_ret_2_0,
      io_ret_2_1 => shiftrows10_io_ret_2_1,
      io_ret_2_2 => shiftrows10_io_ret_2_2,
      io_ret_2_3 => shiftrows10_io_ret_2_3,
      io_ret_3_0 => shiftrows10_io_ret_3_0,
      io_ret_3_1 => shiftrows10_io_ret_3_1,
      io_ret_3_2 => shiftrows10_io_ret_3_2,
      io_ret_3_3 => shiftrows10_io_ret_3_3 
    );
  addroundkey10 : entity work.AddRoundKey
    port map ( 
      io_rk_0_0 => keyschedule9_io_ret_0_0,
      io_rk_0_1 => keyschedule9_io_ret_0_1,
      io_rk_0_2 => keyschedule9_io_ret_0_2,
      io_rk_0_3 => keyschedule9_io_ret_0_3,
      io_rk_1_0 => keyschedule9_io_ret_1_0,
      io_rk_1_1 => keyschedule9_io_ret_1_1,
      io_rk_1_2 => keyschedule9_io_ret_1_2,
      io_rk_1_3 => keyschedule9_io_ret_1_3,
      io_rk_2_0 => keyschedule9_io_ret_2_0,
      io_rk_2_1 => keyschedule9_io_ret_2_1,
      io_rk_2_2 => keyschedule9_io_ret_2_2,
      io_rk_2_3 => keyschedule9_io_ret_2_3,
      io_rk_3_0 => keyschedule9_io_ret_3_0,
      io_rk_3_1 => keyschedule9_io_ret_3_1,
      io_rk_3_2 => keyschedule9_io_ret_3_2,
      io_rk_3_3 => keyschedule9_io_ret_3_3,
      io_s_0_0 => shiftrows10_io_ret_0_0,
      io_s_0_1 => shiftrows10_io_ret_0_1,
      io_s_0_2 => shiftrows10_io_ret_0_2,
      io_s_0_3 => shiftrows10_io_ret_0_3,
      io_s_1_0 => shiftrows10_io_ret_1_0,
      io_s_1_1 => shiftrows10_io_ret_1_1,
      io_s_1_2 => shiftrows10_io_ret_1_2,
      io_s_1_3 => shiftrows10_io_ret_1_3,
      io_s_2_0 => shiftrows10_io_ret_2_0,
      io_s_2_1 => shiftrows10_io_ret_2_1,
      io_s_2_2 => shiftrows10_io_ret_2_2,
      io_s_2_3 => shiftrows10_io_ret_2_3,
      io_s_3_0 => shiftrows10_io_ret_3_0,
      io_s_3_1 => shiftrows10_io_ret_3_1,
      io_s_3_2 => shiftrows10_io_ret_3_2,
      io_s_3_3 => shiftrows10_io_ret_3_3,
      io_ret_0_0 => addroundkey10_io_ret_0_0,
      io_ret_0_1 => addroundkey10_io_ret_0_1,
      io_ret_0_2 => addroundkey10_io_ret_0_2,
      io_ret_0_3 => addroundkey10_io_ret_0_3,
      io_ret_1_0 => addroundkey10_io_ret_1_0,
      io_ret_1_1 => addroundkey10_io_ret_1_1,
      io_ret_1_2 => addroundkey10_io_ret_1_2,
      io_ret_1_3 => addroundkey10_io_ret_1_3,
      io_ret_2_0 => addroundkey10_io_ret_2_0,
      io_ret_2_1 => addroundkey10_io_ret_2_1,
      io_ret_2_2 => addroundkey10_io_ret_2_2,
      io_ret_2_3 => addroundkey10_io_ret_2_3,
      io_ret_3_0 => addroundkey10_io_ret_3_0,
      io_ret_3_1 => addroundkey10_io_ret_3_1,
      io_ret_3_2 => addroundkey10_io_ret_3_2,
      io_ret_3_3 => addroundkey10_io_ret_3_3 
    );
  rcs0 <= pkg_stdLogicVector("00000001");
  keys0_0_0 <= pkg_extract(io_key,127,120);
  keys0_0_1 <= pkg_extract(io_key,95,88);
  keys0_0_2 <= pkg_extract(io_key,63,56);
  keys0_0_3 <= pkg_extract(io_key,31,24);
  keys0_1_0 <= pkg_extract(io_key,119,112);
  keys0_1_1 <= pkg_extract(io_key,87,80);
  keys0_1_2 <= pkg_extract(io_key,55,48);
  keys0_1_3 <= pkg_extract(io_key,23,16);
  keys0_2_0 <= pkg_extract(io_key,111,104);
  keys0_2_1 <= pkg_extract(io_key,79,72);
  keys0_2_2 <= pkg_extract(io_key,47,40);
  keys0_2_3 <= pkg_extract(io_key,15,8);
  keys0_3_0 <= pkg_extract(io_key,103,96);
  keys0_3_1 <= pkg_extract(io_key,71,64);
  keys0_3_2 <= pkg_extract(io_key,39,32);
  keys0_3_3 <= pkg_extract(io_key,7,0);
  addroundkey0_io_s_0_0 <= pkg_extract(io_pt,127,120);
  addroundkey0_io_s_0_1 <= pkg_extract(io_pt,95,88);
  addroundkey0_io_s_0_2 <= pkg_extract(io_pt,63,56);
  addroundkey0_io_s_0_3 <= pkg_extract(io_pt,31,24);
  addroundkey0_io_s_1_0 <= pkg_extract(io_pt,119,112);
  addroundkey0_io_s_1_1 <= pkg_extract(io_pt,87,80);
  addroundkey0_io_s_1_2 <= pkg_extract(io_pt,55,48);
  addroundkey0_io_s_1_3 <= pkg_extract(io_pt,23,16);
  addroundkey0_io_s_2_0 <= pkg_extract(io_pt,111,104);
  addroundkey0_io_s_2_1 <= pkg_extract(io_pt,79,72);
  addroundkey0_io_s_2_2 <= pkg_extract(io_pt,47,40);
  addroundkey0_io_s_2_3 <= pkg_extract(io_pt,15,8);
  addroundkey0_io_s_3_0 <= pkg_extract(io_pt,103,96);
  addroundkey0_io_s_3_1 <= pkg_extract(io_pt,71,64);
  addroundkey0_io_s_3_2 <= pkg_extract(io_pt,39,32);
  addroundkey0_io_s_3_3 <= pkg_extract(io_pt,7,0);
  state0_0_0 <= addroundkey0_io_ret_0_0;
  state0_0_1 <= addroundkey0_io_ret_0_1;
  state0_0_2 <= addroundkey0_io_ret_0_2;
  state0_0_3 <= addroundkey0_io_ret_0_3;
  state0_1_0 <= addroundkey0_io_ret_1_0;
  state0_1_1 <= addroundkey0_io_ret_1_1;
  state0_1_2 <= addroundkey0_io_ret_1_2;
  state0_1_3 <= addroundkey0_io_ret_1_3;
  state0_2_0 <= addroundkey0_io_ret_2_0;
  state0_2_1 <= addroundkey0_io_ret_2_1;
  state0_2_2 <= addroundkey0_io_ret_2_2;
  state0_2_3 <= addroundkey0_io_ret_2_3;
  state0_3_0 <= addroundkey0_io_ret_3_0;
  state0_3_1 <= addroundkey0_io_ret_3_1;
  state0_3_2 <= addroundkey0_io_ret_3_2;
  state0_3_3 <= addroundkey0_io_ret_3_3;
  process(addroundkey10_io_ret_0_0,addroundkey10_io_ret_0_1,addroundkey10_io_ret_0_2,addroundkey10_io_ret_0_3,addroundkey10_io_ret_1_0,addroundkey10_io_ret_1_1,addroundkey10_io_ret_1_2,addroundkey10_io_ret_1_3,addroundkey10_io_ret_2_0,addroundkey10_io_ret_2_1,addroundkey10_io_ret_2_2,addroundkey10_io_ret_2_3,addroundkey10_io_ret_3_0,addroundkey10_io_ret_3_1,addroundkey10_io_ret_3_2,addroundkey10_io_ret_3_3)
  begin
    zz_io_ret(127 downto 120) <= addroundkey10_io_ret_0_0;
    zz_io_ret(95 downto 88) <= addroundkey10_io_ret_0_1;
    zz_io_ret(63 downto 56) <= addroundkey10_io_ret_0_2;
    zz_io_ret(31 downto 24) <= addroundkey10_io_ret_0_3;
    zz_io_ret(119 downto 112) <= addroundkey10_io_ret_1_0;
    zz_io_ret(87 downto 80) <= addroundkey10_io_ret_1_1;
    zz_io_ret(55 downto 48) <= addroundkey10_io_ret_1_2;
    zz_io_ret(23 downto 16) <= addroundkey10_io_ret_1_3;
    zz_io_ret(111 downto 104) <= addroundkey10_io_ret_2_0;
    zz_io_ret(79 downto 72) <= addroundkey10_io_ret_2_1;
    zz_io_ret(47 downto 40) <= addroundkey10_io_ret_2_2;
    zz_io_ret(15 downto 8) <= addroundkey10_io_ret_2_3;
    zz_io_ret(103 downto 96) <= addroundkey10_io_ret_3_0;
    zz_io_ret(71 downto 64) <= addroundkey10_io_ret_3_1;
    zz_io_ret(39 downto 32) <= addroundkey10_io_ret_3_2;
    zz_io_ret(7 downto 0) <= addroundkey10_io_ret_3_3;
  end process;

  io_ret <= zz_io_ret;
end arch;

