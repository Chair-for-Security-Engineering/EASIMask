-- Generator : SpinalHDL v1.6.2    git head : e20135930d099f5d7469bbea4f2ca5d14698f642
-- Component : G256InvTIMaskedN
-- Git hash  : e20135930d099f5d7469bbea4f2ca5d14698f642

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;

package pkg_enum is

end pkg_enum;

library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

package pkg_scala2hdl is
  function pkg_extract (that : std_logic_vector; bitId : integer) return std_logic;
  function pkg_extract (that : std_logic_vector; base : unsigned; size : integer) return std_logic_vector;
  function pkg_cat (a : std_logic_vector; b : std_logic_vector) return std_logic_vector;
  function pkg_not (value : std_logic_vector) return std_logic_vector;
  function pkg_extract (that : unsigned; bitId : integer) return std_logic;
  function pkg_extract (that : unsigned; base : unsigned; size : integer) return unsigned;
  function pkg_cat (a : unsigned; b : unsigned) return unsigned;
  function pkg_not (value : unsigned) return unsigned;
  function pkg_extract (that : signed; bitId : integer) return std_logic;
  function pkg_extract (that : signed; base : unsigned; size : integer) return signed;
  function pkg_cat (a : signed; b : signed) return signed;
  function pkg_not (value : signed) return signed;

  function pkg_mux (sel : std_logic; one : std_logic; zero : std_logic) return std_logic;
  function pkg_mux (sel : std_logic; one : std_logic_vector; zero : std_logic_vector) return std_logic_vector;
  function pkg_mux (sel : std_logic; one : unsigned; zero : unsigned) return unsigned;
  function pkg_mux (sel : std_logic; one : signed; zero : signed) return signed;

  function pkg_toStdLogic (value : boolean) return std_logic;
  function pkg_toStdLogicVector (value : std_logic) return std_logic_vector;
  function pkg_toUnsigned (value : std_logic) return unsigned;
  function pkg_toSigned (value : std_logic) return signed;
  function pkg_stdLogicVector (lit : std_logic_vector) return std_logic_vector;
  function pkg_unsigned (lit : unsigned) return unsigned;
  function pkg_signed (lit : signed) return signed;

  function pkg_resize (that : std_logic_vector; width : integer) return std_logic_vector;
  function pkg_resize (that : unsigned; width : integer) return unsigned;
  function pkg_resize (that : signed; width : integer) return signed;

  function pkg_extract (that : std_logic_vector; high : integer; low : integer) return std_logic_vector;
  function pkg_extract (that : unsigned; high : integer; low : integer) return unsigned;
  function pkg_extract (that : signed; high : integer; low : integer) return signed;

  function pkg_shiftRight (that : std_logic_vector; size : natural) return std_logic_vector;
  function pkg_shiftRight (that : std_logic_vector; size : unsigned) return std_logic_vector;
  function pkg_shiftLeft (that : std_logic_vector; size : natural) return std_logic_vector;
  function pkg_shiftLeft (that : std_logic_vector; size : unsigned) return std_logic_vector;

  function pkg_shiftRight (that : unsigned; size : natural) return unsigned;
  function pkg_shiftRight (that : unsigned; size : unsigned) return unsigned;
  function pkg_shiftLeft (that : unsigned; size : natural) return unsigned;
  function pkg_shiftLeft (that : unsigned; size : unsigned) return unsigned;

  function pkg_shiftRight (that : signed; size : natural) return signed;
  function pkg_shiftRight (that : signed; size : unsigned) return signed;
  function pkg_shiftLeft (that : signed; size : natural) return signed;
  function pkg_shiftLeft (that : signed; size : unsigned; w : integer) return signed;

  function pkg_rotateLeft (that : std_logic_vector; size : unsigned) return std_logic_vector;
end  pkg_scala2hdl;

package body pkg_scala2hdl is
  function pkg_extract (that : std_logic_vector; bitId : integer) return std_logic is
    alias temp : std_logic_vector(that'length-1 downto 0) is that;
  begin
    return temp(bitId);
  end pkg_extract;

  function pkg_extract (that : std_logic_vector; base : unsigned; size : integer) return std_logic_vector is
    alias temp : std_logic_vector(that'length-1 downto 0) is that;    constant elementCount : integer := temp'length - size + 1;
    type tableType is array (0 to elementCount-1) of std_logic_vector(size-1 downto 0);
    variable table : tableType;
  begin
    for i in 0 to elementCount-1 loop
      table(i) := temp(i + size - 1 downto i);
    end loop;
    return table(to_integer(base));
  end pkg_extract;

  function pkg_cat (a : std_logic_vector; b : std_logic_vector) return std_logic_vector is
    variable cat : std_logic_vector(a'length + b'length-1 downto 0);
  begin
    cat := a & b;
    return cat;
  end pkg_cat;

  function pkg_not (value : std_logic_vector) return std_logic_vector is
    variable ret : std_logic_vector(value'length-1 downto 0);
  begin
    ret := not value;
    return ret;
  end pkg_not;

  function pkg_extract (that : unsigned; bitId : integer) return std_logic is
    alias temp : unsigned(that'length-1 downto 0) is that;
  begin
    return temp(bitId);
  end pkg_extract;

  function pkg_extract (that : unsigned; base : unsigned; size : integer) return unsigned is
    alias temp : unsigned(that'length-1 downto 0) is that;    constant elementCount : integer := temp'length - size + 1;
    type tableType is array (0 to elementCount-1) of unsigned(size-1 downto 0);
    variable table : tableType;
  begin
    for i in 0 to elementCount-1 loop
      table(i) := temp(i + size - 1 downto i);
    end loop;
    return table(to_integer(base));
  end pkg_extract;

  function pkg_cat (a : unsigned; b : unsigned) return unsigned is
    variable cat : unsigned(a'length + b'length-1 downto 0);
  begin
    cat := a & b;
    return cat;
  end pkg_cat;

  function pkg_not (value : unsigned) return unsigned is
    variable ret : unsigned(value'length-1 downto 0);
  begin
    ret := not value;
    return ret;
  end pkg_not;

  function pkg_extract (that : signed; bitId : integer) return std_logic is
    alias temp : signed(that'length-1 downto 0) is that;
  begin
    return temp(bitId);
  end pkg_extract;

  function pkg_extract (that : signed; base : unsigned; size : integer) return signed is
    alias temp : signed(that'length-1 downto 0) is that;    constant elementCount : integer := temp'length - size + 1;
    type tableType is array (0 to elementCount-1) of signed(size-1 downto 0);
    variable table : tableType;
  begin
    for i in 0 to elementCount-1 loop
      table(i) := temp(i + size - 1 downto i);
    end loop;
    return table(to_integer(base));
  end pkg_extract;

  function pkg_cat (a : signed; b : signed) return signed is
    variable cat : signed(a'length + b'length-1 downto 0);
  begin
    cat := a & b;
    return cat;
  end pkg_cat;

  function pkg_not (value : signed) return signed is
    variable ret : signed(value'length-1 downto 0);
  begin
    ret := not value;
    return ret;
  end pkg_not;


  -- unsigned shifts
  function pkg_shiftRight (that : unsigned; size : natural) return unsigned is
    variable ret : unsigned(that'length-1 downto 0);
  begin
    if size >= that'length then
      return "";
    else
      ret := shift_right(that,size);
      return ret(that'length-1-size downto 0);
    end if;
  end pkg_shiftRight;

  function pkg_shiftRight (that : unsigned; size : unsigned) return unsigned is
    variable ret : unsigned(that'length-1 downto 0);
  begin
    ret := shift_right(that,to_integer(size));
    return ret;
  end pkg_shiftRight;

  function pkg_shiftLeft (that : unsigned; size : natural) return unsigned is
  begin
    return shift_left(resize(that,that'length + size),size);
  end pkg_shiftLeft;

  function pkg_shiftLeft (that : unsigned; size : unsigned) return unsigned is
  begin
    return shift_left(resize(that,that'length + 2**size'length - 1),to_integer(size));
  end pkg_shiftLeft;

  -- std_logic_vector shifts
  function pkg_shiftRight (that : std_logic_vector; size : natural) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftRight(unsigned(that),size));
  end pkg_shiftRight;

  function pkg_shiftRight (that : std_logic_vector; size : unsigned) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftRight(unsigned(that),size));
  end pkg_shiftRight;

  function pkg_shiftLeft (that : std_logic_vector; size : natural) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftLeft(unsigned(that),size));
  end pkg_shiftLeft;

  function pkg_shiftLeft (that : std_logic_vector; size : unsigned) return std_logic_vector is
  begin
    return std_logic_vector(pkg_shiftLeft(unsigned(that),size));
  end pkg_shiftLeft;

  -- signed shifts
  function pkg_shiftRight (that : signed; size : natural) return signed is
  begin
    return signed(pkg_shiftRight(unsigned(that),size));
  end pkg_shiftRight;

  function pkg_shiftRight (that : signed; size : unsigned) return signed is
  begin
    return shift_right(that,to_integer(size));
  end pkg_shiftRight;

  function pkg_shiftLeft (that : signed; size : natural) return signed is
  begin
    return signed(pkg_shiftLeft(unsigned(that),size));
  end pkg_shiftLeft;

  function pkg_shiftLeft (that : signed; size : unsigned; w : integer) return signed is
  begin
    return shift_left(resize(that,w),to_integer(size));
  end pkg_shiftLeft;

  function pkg_rotateLeft (that : std_logic_vector; size : unsigned) return std_logic_vector is
  begin
    return std_logic_vector(rotate_left(unsigned(that),to_integer(size)));
  end pkg_rotateLeft;

  function pkg_extract (that : std_logic_vector; high : integer; low : integer) return std_logic_vector is
    alias temp : std_logic_vector(that'length-1 downto 0) is that;
  begin
    return temp(high downto low);
  end pkg_extract;

  function pkg_extract (that : unsigned; high : integer; low : integer) return unsigned is
    alias temp : unsigned(that'length-1 downto 0) is that;
  begin
    return temp(high downto low);
  end pkg_extract;

  function pkg_extract (that : signed; high : integer; low : integer) return signed is
    alias temp : signed(that'length-1 downto 0) is that;
  begin
    return temp(high downto low);
  end pkg_extract;

  function pkg_mux (sel : std_logic; one : std_logic; zero : std_logic) return std_logic is
  begin
    if sel = '1' then
      return one;
    else
      return zero;
    end if;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : std_logic_vector; zero : std_logic_vector) return std_logic_vector is
    variable ret : std_logic_vector(zero'range);
  begin
    if sel = '1' then
      ret := one;
    else
      ret := zero;
    end if;
    return ret;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : unsigned; zero : unsigned) return unsigned is
    variable ret : unsigned(zero'range);
  begin
    if sel = '1' then
      ret := one;
    else
      ret := zero;
    end if;
    return ret;
  end pkg_mux;

  function pkg_mux (sel : std_logic; one : signed; zero : signed) return signed is
    variable ret : signed(zero'range);
  begin
    if sel = '1' then
      ret := one;
    else
      ret := zero;
    end if;
    return ret;
  end pkg_mux;

  function pkg_toStdLogic (value : boolean) return std_logic is
  begin
    if value = true then
      return '1';
    else
      return '0';
    end if;
  end pkg_toStdLogic;

  function pkg_toStdLogicVector (value : std_logic) return std_logic_vector is
    variable ret : std_logic_vector(0 downto 0);
  begin
    ret(0) := value;
    return ret;
  end pkg_toStdLogicVector;

  function pkg_toUnsigned (value : std_logic) return unsigned is
    variable ret : unsigned(0 downto 0);
  begin
    ret(0) := value;
    return ret;
  end pkg_toUnsigned;

  function pkg_toSigned (value : std_logic) return signed is
    variable ret : signed(0 downto 0);
  begin
    ret(0) := value;
    return ret;
  end pkg_toSigned;

  function pkg_stdLogicVector (lit : std_logic_vector) return std_logic_vector is
    alias ret : std_logic_vector(lit'length-1 downto 0) is lit;
  begin
    return ret;
  end pkg_stdLogicVector;

  function pkg_unsigned (lit : unsigned) return unsigned is
    alias ret : unsigned(lit'length-1 downto 0) is lit;
  begin
    return ret;
  end pkg_unsigned;

  function pkg_signed (lit : signed) return signed is
    alias ret : signed(lit'length-1 downto 0) is lit;
  begin
    return ret;
  end pkg_signed;

  function pkg_resize (that : std_logic_vector; width : integer) return std_logic_vector is
  begin
    return std_logic_vector(resize(unsigned(that),width));
  end pkg_resize;

  function pkg_resize (that : unsigned; width : integer) return unsigned is
    variable ret : unsigned(width-1 downto 0);
  begin
    if that'length = 0 then
       ret := (others => '0');
    else
       ret := resize(that,width);
    end if;
    return ret;
  end pkg_resize;
  function pkg_resize (that : signed; width : integer) return signed is
    alias temp : signed(that'length-1 downto 0) is that;
    variable ret : signed(width-1 downto 0);
  begin
    if temp'length = 0 then
       ret := (others => '0');
    elsif temp'length >= width then
       ret := temp(width-1 downto 0);
    else
       ret := resize(temp,width);
    end if;
    return ret;
  end pkg_resize;
end pkg_scala2hdl;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity G4MulTIMaskedN is
  port(
    io_x_0 : in std_logic_vector(1 downto 0);
    io_x_1 : in std_logic_vector(1 downto 0);
    io_x_2 : in std_logic_vector(1 downto 0);
    io_x_3 : in std_logic_vector(1 downto 0);
    io_x_4 : in std_logic_vector(1 downto 0);
    io_x_5 : in std_logic_vector(1 downto 0);
    io_x_6 : in std_logic_vector(1 downto 0);
    io_x_7 : in std_logic_vector(1 downto 0);
    io_x_8 : in std_logic_vector(1 downto 0);
    io_x_9 : in std_logic_vector(1 downto 0);
    io_x_10 : in std_logic_vector(1 downto 0);
    io_x_11 : in std_logic_vector(1 downto 0);
    io_x_12 : in std_logic_vector(1 downto 0);
    io_y_0 : in std_logic_vector(1 downto 0);
    io_y_1 : in std_logic_vector(1 downto 0);
    io_y_2 : in std_logic_vector(1 downto 0);
    io_y_3 : in std_logic_vector(1 downto 0);
    io_y_4 : in std_logic_vector(1 downto 0);
    io_y_5 : in std_logic_vector(1 downto 0);
    io_y_6 : in std_logic_vector(1 downto 0);
    io_y_7 : in std_logic_vector(1 downto 0);
    io_y_8 : in std_logic_vector(1 downto 0);
    io_y_9 : in std_logic_vector(1 downto 0);
    io_y_10 : in std_logic_vector(1 downto 0);
    io_y_11 : in std_logic_vector(1 downto 0);
    io_y_12 : in std_logic_vector(1 downto 0);
    io_z_0 : out std_logic_vector(1 downto 0);
    io_z_1 : out std_logic_vector(1 downto 0);
    io_z_2 : out std_logic_vector(1 downto 0);
    io_z_3 : out std_logic_vector(1 downto 0);
    io_z_4 : out std_logic_vector(1 downto 0);
    io_z_5 : out std_logic_vector(1 downto 0);
    io_z_6 : out std_logic_vector(1 downto 0);
    io_z_7 : out std_logic_vector(1 downto 0);
    io_z_8 : out std_logic_vector(1 downto 0);
    io_z_9 : out std_logic_vector(1 downto 0);
    io_z_10 : out std_logic_vector(1 downto 0);
    io_z_11 : out std_logic_vector(1 downto 0);
    io_z_12 : out std_logic_vector(1 downto 0);
    clk : in std_logic;
    reset : in std_logic
  );
end G4MulTIMaskedN;

architecture arch of G4MulTIMaskedN is

  signal dummy : std_logic;
  signal a_0 : std_logic;
  signal a_1 : std_logic;
  signal a_2 : std_logic;
  signal a_3 : std_logic;
  signal a_4 : std_logic;
  signal a_5 : std_logic;
  signal a_6 : std_logic;
  signal a_7 : std_logic;
  signal a_8 : std_logic;
  signal a_9 : std_logic;
  signal a_10 : std_logic;
  signal a_11 : std_logic;
  signal a_12 : std_logic;
  signal b_0 : std_logic;
  signal b_1 : std_logic;
  signal b_2 : std_logic;
  signal b_3 : std_logic;
  signal b_4 : std_logic;
  signal b_5 : std_logic;
  signal b_6 : std_logic;
  signal b_7 : std_logic;
  signal b_8 : std_logic;
  signal b_9 : std_logic;
  signal b_10 : std_logic;
  signal b_11 : std_logic;
  signal b_12 : std_logic;
  signal c_0 : std_logic;
  signal c_1 : std_logic;
  signal c_2 : std_logic;
  signal c_3 : std_logic;
  signal c_4 : std_logic;
  signal c_5 : std_logic;
  signal c_6 : std_logic;
  signal c_7 : std_logic;
  signal c_8 : std_logic;
  signal c_9 : std_logic;
  signal c_10 : std_logic;
  signal c_11 : std_logic;
  signal c_12 : std_logic;
  signal d_0 : std_logic;
  signal d_1 : std_logic;
  signal d_2 : std_logic;
  signal d_3 : std_logic;
  signal d_4 : std_logic;
  signal d_5 : std_logic;
  signal d_6 : std_logic;
  signal d_7 : std_logic;
  signal d_8 : std_logic;
  signal d_9 : std_logic;
  signal d_10 : std_logic;
  signal d_11 : std_logic;
  signal d_12 : std_logic;
  signal e_0 : std_logic_vector(12 downto 0);
  signal e_1 : std_logic_vector(12 downto 0);
  signal e_2 : std_logic_vector(12 downto 0);
  signal e_3 : std_logic_vector(12 downto 0);
  signal e_4 : std_logic_vector(12 downto 0);
  signal e_5 : std_logic_vector(12 downto 0);
  signal e_6 : std_logic_vector(12 downto 0);
  signal e_7 : std_logic_vector(12 downto 0);
  signal e_8 : std_logic_vector(12 downto 0);
  signal e_9 : std_logic_vector(12 downto 0);
  signal e_10 : std_logic_vector(12 downto 0);
  signal e_11 : std_logic_vector(12 downto 0);
  signal e_12 : std_logic_vector(12 downto 0);
  signal f_0 : std_logic_vector(12 downto 0);
  signal f_1 : std_logic_vector(12 downto 0);
  signal f_2 : std_logic_vector(12 downto 0);
  signal f_3 : std_logic_vector(12 downto 0);
  signal f_4 : std_logic_vector(12 downto 0);
  signal f_5 : std_logic_vector(12 downto 0);
  signal f_6 : std_logic_vector(12 downto 0);
  signal f_7 : std_logic_vector(12 downto 0);
  signal f_8 : std_logic_vector(12 downto 0);
  signal f_9 : std_logic_vector(12 downto 0);
  signal f_10 : std_logic_vector(12 downto 0);
  signal f_11 : std_logic_vector(12 downto 0);
  signal f_12 : std_logic_vector(12 downto 0);
  signal ac_0 : std_logic;
  signal ac_1 : std_logic;
  signal ac_2 : std_logic;
  signal ac_3 : std_logic;
  signal ac_4 : std_logic;
  signal ac_5 : std_logic;
  signal ac_6 : std_logic;
  signal ac_7 : std_logic;
  signal ac_8 : std_logic;
  signal ac_9 : std_logic;
  signal ac_10 : std_logic;
  signal ac_11 : std_logic;
  signal ac_12 : std_logic;
  signal ac_13 : std_logic;
  signal ac_14 : std_logic;
  signal ac_15 : std_logic;
  signal ac_16 : std_logic;
  signal ac_17 : std_logic;
  signal ac_18 : std_logic;
  signal ac_19 : std_logic;
  signal ac_20 : std_logic;
  signal ac_21 : std_logic;
  signal ac_22 : std_logic;
  signal ac_23 : std_logic;
  signal ac_24 : std_logic;
  signal ac_25 : std_logic;
  signal ac_26 : std_logic;
  signal ac_27 : std_logic;
  signal ac_28 : std_logic;
  signal ac_29 : std_logic;
  signal ac_30 : std_logic;
  signal ac_31 : std_logic;
  signal ac_32 : std_logic;
  signal ac_33 : std_logic;
  signal ac_34 : std_logic;
  signal ac_35 : std_logic;
  signal ac_36 : std_logic;
  signal ac_37 : std_logic;
  signal ac_38 : std_logic;
  signal ac_39 : std_logic;
  signal ac_40 : std_logic;
  signal ac_41 : std_logic;
  signal ac_42 : std_logic;
  signal ac_43 : std_logic;
  signal ac_44 : std_logic;
  signal ac_45 : std_logic;
  signal ac_46 : std_logic;
  signal ac_47 : std_logic;
  signal ac_48 : std_logic;
  signal ac_49 : std_logic;
  signal ac_50 : std_logic;
  signal ac_51 : std_logic;
  signal ac_52 : std_logic;
  signal ac_53 : std_logic;
  signal ac_54 : std_logic;
  signal ac_55 : std_logic;
  signal ac_56 : std_logic;
  signal ac_57 : std_logic;
  signal ac_58 : std_logic;
  signal ac_59 : std_logic;
  signal ac_60 : std_logic;
  signal ac_61 : std_logic;
  signal ac_62 : std_logic;
  signal ac_63 : std_logic;
  signal ac_64 : std_logic;
  signal ac_65 : std_logic;
  signal ac_66 : std_logic;
  signal ac_67 : std_logic;
  signal ac_68 : std_logic;
  signal ac_69 : std_logic;
  signal ac_70 : std_logic;
  signal ac_71 : std_logic;
  signal ac_72 : std_logic;
  signal ac_73 : std_logic;
  signal ac_74 : std_logic;
  signal ac_75 : std_logic;
  signal ac_76 : std_logic;
  signal ac_77 : std_logic;
  signal ac_78 : std_logic;
  signal ac_79 : std_logic;
  signal ac_80 : std_logic;
  signal ac_81 : std_logic;
  signal ac_82 : std_logic;
  signal ac_83 : std_logic;
  signal ac_84 : std_logic;
  signal ac_85 : std_logic;
  signal ac_86 : std_logic;
  signal ac_87 : std_logic;
  signal ac_88 : std_logic;
  signal ac_89 : std_logic;
  signal ac_90 : std_logic;
  signal ac_91 : std_logic;
  signal ac_92 : std_logic;
  signal ac_93 : std_logic;
  signal ac_94 : std_logic;
  signal ac_95 : std_logic;
  signal ac_96 : std_logic;
  signal ac_97 : std_logic;
  signal ac_98 : std_logic;
  signal ac_99 : std_logic;
  signal ac_100 : std_logic;
  signal ac_101 : std_logic;
  signal ac_102 : std_logic;
  signal ac_103 : std_logic;
  signal ac_104 : std_logic;
  signal ac_105 : std_logic;
  signal ac_106 : std_logic;
  signal ac_107 : std_logic;
  signal ac_108 : std_logic;
  signal ac_109 : std_logic;
  signal ac_110 : std_logic;
  signal ac_111 : std_logic;
  signal ac_112 : std_logic;
  signal ac_113 : std_logic;
  signal ac_114 : std_logic;
  signal ac_115 : std_logic;
  signal ac_116 : std_logic;
  signal ac_117 : std_logic;
  signal ac_118 : std_logic;
  signal ac_119 : std_logic;
  signal ac_120 : std_logic;
  signal ac_121 : std_logic;
  signal ac_122 : std_logic;
  signal ac_123 : std_logic;
  signal ac_124 : std_logic;
  signal ac_125 : std_logic;
  signal ac_126 : std_logic;
  signal ac_127 : std_logic;
  signal ac_128 : std_logic;
  signal ac_129 : std_logic;
  signal ac_130 : std_logic;
  signal ac_131 : std_logic;
  signal ac_132 : std_logic;
  signal ac_133 : std_logic;
  signal ac_134 : std_logic;
  signal ac_135 : std_logic;
  signal ac_136 : std_logic;
  signal ac_137 : std_logic;
  signal ac_138 : std_logic;
  signal ac_139 : std_logic;
  signal ac_140 : std_logic;
  signal ac_141 : std_logic;
  signal ac_142 : std_logic;
  signal ac_143 : std_logic;
  signal ac_144 : std_logic;
  signal ac_145 : std_logic;
  signal ac_146 : std_logic;
  signal ac_147 : std_logic;
  signal ac_148 : std_logic;
  signal ac_149 : std_logic;
  signal ac_150 : std_logic;
  signal ac_151 : std_logic;
  signal ac_152 : std_logic;
  signal ac_153 : std_logic;
  signal ac_154 : std_logic;
  signal ac_155 : std_logic;
  signal ac_156 : std_logic;
  signal ac_157 : std_logic;
  signal ac_158 : std_logic;
  signal ac_159 : std_logic;
  signal ac_160 : std_logic;
  signal ac_161 : std_logic;
  signal ac_162 : std_logic;
  signal ac_163 : std_logic;
  signal ac_164 : std_logic;
  signal ac_165 : std_logic;
  signal ac_166 : std_logic;
  signal ac_167 : std_logic;
  signal ac_168 : std_logic;
  signal ad_0 : std_logic;
  signal ad_1 : std_logic;
  signal ad_2 : std_logic;
  signal ad_3 : std_logic;
  signal ad_4 : std_logic;
  signal ad_5 : std_logic;
  signal ad_6 : std_logic;
  signal ad_7 : std_logic;
  signal ad_8 : std_logic;
  signal ad_9 : std_logic;
  signal ad_10 : std_logic;
  signal ad_11 : std_logic;
  signal ad_12 : std_logic;
  signal ad_13 : std_logic;
  signal ad_14 : std_logic;
  signal ad_15 : std_logic;
  signal ad_16 : std_logic;
  signal ad_17 : std_logic;
  signal ad_18 : std_logic;
  signal ad_19 : std_logic;
  signal ad_20 : std_logic;
  signal ad_21 : std_logic;
  signal ad_22 : std_logic;
  signal ad_23 : std_logic;
  signal ad_24 : std_logic;
  signal ad_25 : std_logic;
  signal ad_26 : std_logic;
  signal ad_27 : std_logic;
  signal ad_28 : std_logic;
  signal ad_29 : std_logic;
  signal ad_30 : std_logic;
  signal ad_31 : std_logic;
  signal ad_32 : std_logic;
  signal ad_33 : std_logic;
  signal ad_34 : std_logic;
  signal ad_35 : std_logic;
  signal ad_36 : std_logic;
  signal ad_37 : std_logic;
  signal ad_38 : std_logic;
  signal ad_39 : std_logic;
  signal ad_40 : std_logic;
  signal ad_41 : std_logic;
  signal ad_42 : std_logic;
  signal ad_43 : std_logic;
  signal ad_44 : std_logic;
  signal ad_45 : std_logic;
  signal ad_46 : std_logic;
  signal ad_47 : std_logic;
  signal ad_48 : std_logic;
  signal ad_49 : std_logic;
  signal ad_50 : std_logic;
  signal ad_51 : std_logic;
  signal ad_52 : std_logic;
  signal ad_53 : std_logic;
  signal ad_54 : std_logic;
  signal ad_55 : std_logic;
  signal ad_56 : std_logic;
  signal ad_57 : std_logic;
  signal ad_58 : std_logic;
  signal ad_59 : std_logic;
  signal ad_60 : std_logic;
  signal ad_61 : std_logic;
  signal ad_62 : std_logic;
  signal ad_63 : std_logic;
  signal ad_64 : std_logic;
  signal ad_65 : std_logic;
  signal ad_66 : std_logic;
  signal ad_67 : std_logic;
  signal ad_68 : std_logic;
  signal ad_69 : std_logic;
  signal ad_70 : std_logic;
  signal ad_71 : std_logic;
  signal ad_72 : std_logic;
  signal ad_73 : std_logic;
  signal ad_74 : std_logic;
  signal ad_75 : std_logic;
  signal ad_76 : std_logic;
  signal ad_77 : std_logic;
  signal ad_78 : std_logic;
  signal ad_79 : std_logic;
  signal ad_80 : std_logic;
  signal ad_81 : std_logic;
  signal ad_82 : std_logic;
  signal ad_83 : std_logic;
  signal ad_84 : std_logic;
  signal ad_85 : std_logic;
  signal ad_86 : std_logic;
  signal ad_87 : std_logic;
  signal ad_88 : std_logic;
  signal ad_89 : std_logic;
  signal ad_90 : std_logic;
  signal ad_91 : std_logic;
  signal ad_92 : std_logic;
  signal ad_93 : std_logic;
  signal ad_94 : std_logic;
  signal ad_95 : std_logic;
  signal ad_96 : std_logic;
  signal ad_97 : std_logic;
  signal ad_98 : std_logic;
  signal ad_99 : std_logic;
  signal ad_100 : std_logic;
  signal ad_101 : std_logic;
  signal ad_102 : std_logic;
  signal ad_103 : std_logic;
  signal ad_104 : std_logic;
  signal ad_105 : std_logic;
  signal ad_106 : std_logic;
  signal ad_107 : std_logic;
  signal ad_108 : std_logic;
  signal ad_109 : std_logic;
  signal ad_110 : std_logic;
  signal ad_111 : std_logic;
  signal ad_112 : std_logic;
  signal ad_113 : std_logic;
  signal ad_114 : std_logic;
  signal ad_115 : std_logic;
  signal ad_116 : std_logic;
  signal ad_117 : std_logic;
  signal ad_118 : std_logic;
  signal ad_119 : std_logic;
  signal ad_120 : std_logic;
  signal ad_121 : std_logic;
  signal ad_122 : std_logic;
  signal ad_123 : std_logic;
  signal ad_124 : std_logic;
  signal ad_125 : std_logic;
  signal ad_126 : std_logic;
  signal ad_127 : std_logic;
  signal ad_128 : std_logic;
  signal ad_129 : std_logic;
  signal ad_130 : std_logic;
  signal ad_131 : std_logic;
  signal ad_132 : std_logic;
  signal ad_133 : std_logic;
  signal ad_134 : std_logic;
  signal ad_135 : std_logic;
  signal ad_136 : std_logic;
  signal ad_137 : std_logic;
  signal ad_138 : std_logic;
  signal ad_139 : std_logic;
  signal ad_140 : std_logic;
  signal ad_141 : std_logic;
  signal ad_142 : std_logic;
  signal ad_143 : std_logic;
  signal ad_144 : std_logic;
  signal ad_145 : std_logic;
  signal ad_146 : std_logic;
  signal ad_147 : std_logic;
  signal ad_148 : std_logic;
  signal ad_149 : std_logic;
  signal ad_150 : std_logic;
  signal ad_151 : std_logic;
  signal ad_152 : std_logic;
  signal ad_153 : std_logic;
  signal ad_154 : std_logic;
  signal ad_155 : std_logic;
  signal ad_156 : std_logic;
  signal ad_157 : std_logic;
  signal ad_158 : std_logic;
  signal ad_159 : std_logic;
  signal ad_160 : std_logic;
  signal ad_161 : std_logic;
  signal ad_162 : std_logic;
  signal ad_163 : std_logic;
  signal ad_164 : std_logic;
  signal ad_165 : std_logic;
  signal ad_166 : std_logic;
  signal ad_167 : std_logic;
  signal ad_168 : std_logic;
  signal bc_0 : std_logic;
  signal bc_1 : std_logic;
  signal bc_2 : std_logic;
  signal bc_3 : std_logic;
  signal bc_4 : std_logic;
  signal bc_5 : std_logic;
  signal bc_6 : std_logic;
  signal bc_7 : std_logic;
  signal bc_8 : std_logic;
  signal bc_9 : std_logic;
  signal bc_10 : std_logic;
  signal bc_11 : std_logic;
  signal bc_12 : std_logic;
  signal bc_13 : std_logic;
  signal bc_14 : std_logic;
  signal bc_15 : std_logic;
  signal bc_16 : std_logic;
  signal bc_17 : std_logic;
  signal bc_18 : std_logic;
  signal bc_19 : std_logic;
  signal bc_20 : std_logic;
  signal bc_21 : std_logic;
  signal bc_22 : std_logic;
  signal bc_23 : std_logic;
  signal bc_24 : std_logic;
  signal bc_25 : std_logic;
  signal bc_26 : std_logic;
  signal bc_27 : std_logic;
  signal bc_28 : std_logic;
  signal bc_29 : std_logic;
  signal bc_30 : std_logic;
  signal bc_31 : std_logic;
  signal bc_32 : std_logic;
  signal bc_33 : std_logic;
  signal bc_34 : std_logic;
  signal bc_35 : std_logic;
  signal bc_36 : std_logic;
  signal bc_37 : std_logic;
  signal bc_38 : std_logic;
  signal bc_39 : std_logic;
  signal bc_40 : std_logic;
  signal bc_41 : std_logic;
  signal bc_42 : std_logic;
  signal bc_43 : std_logic;
  signal bc_44 : std_logic;
  signal bc_45 : std_logic;
  signal bc_46 : std_logic;
  signal bc_47 : std_logic;
  signal bc_48 : std_logic;
  signal bc_49 : std_logic;
  signal bc_50 : std_logic;
  signal bc_51 : std_logic;
  signal bc_52 : std_logic;
  signal bc_53 : std_logic;
  signal bc_54 : std_logic;
  signal bc_55 : std_logic;
  signal bc_56 : std_logic;
  signal bc_57 : std_logic;
  signal bc_58 : std_logic;
  signal bc_59 : std_logic;
  signal bc_60 : std_logic;
  signal bc_61 : std_logic;
  signal bc_62 : std_logic;
  signal bc_63 : std_logic;
  signal bc_64 : std_logic;
  signal bc_65 : std_logic;
  signal bc_66 : std_logic;
  signal bc_67 : std_logic;
  signal bc_68 : std_logic;
  signal bc_69 : std_logic;
  signal bc_70 : std_logic;
  signal bc_71 : std_logic;
  signal bc_72 : std_logic;
  signal bc_73 : std_logic;
  signal bc_74 : std_logic;
  signal bc_75 : std_logic;
  signal bc_76 : std_logic;
  signal bc_77 : std_logic;
  signal bc_78 : std_logic;
  signal bc_79 : std_logic;
  signal bc_80 : std_logic;
  signal bc_81 : std_logic;
  signal bc_82 : std_logic;
  signal bc_83 : std_logic;
  signal bc_84 : std_logic;
  signal bc_85 : std_logic;
  signal bc_86 : std_logic;
  signal bc_87 : std_logic;
  signal bc_88 : std_logic;
  signal bc_89 : std_logic;
  signal bc_90 : std_logic;
  signal bc_91 : std_logic;
  signal bc_92 : std_logic;
  signal bc_93 : std_logic;
  signal bc_94 : std_logic;
  signal bc_95 : std_logic;
  signal bc_96 : std_logic;
  signal bc_97 : std_logic;
  signal bc_98 : std_logic;
  signal bc_99 : std_logic;
  signal bc_100 : std_logic;
  signal bc_101 : std_logic;
  signal bc_102 : std_logic;
  signal bc_103 : std_logic;
  signal bc_104 : std_logic;
  signal bc_105 : std_logic;
  signal bc_106 : std_logic;
  signal bc_107 : std_logic;
  signal bc_108 : std_logic;
  signal bc_109 : std_logic;
  signal bc_110 : std_logic;
  signal bc_111 : std_logic;
  signal bc_112 : std_logic;
  signal bc_113 : std_logic;
  signal bc_114 : std_logic;
  signal bc_115 : std_logic;
  signal bc_116 : std_logic;
  signal bc_117 : std_logic;
  signal bc_118 : std_logic;
  signal bc_119 : std_logic;
  signal bc_120 : std_logic;
  signal bc_121 : std_logic;
  signal bc_122 : std_logic;
  signal bc_123 : std_logic;
  signal bc_124 : std_logic;
  signal bc_125 : std_logic;
  signal bc_126 : std_logic;
  signal bc_127 : std_logic;
  signal bc_128 : std_logic;
  signal bc_129 : std_logic;
  signal bc_130 : std_logic;
  signal bc_131 : std_logic;
  signal bc_132 : std_logic;
  signal bc_133 : std_logic;
  signal bc_134 : std_logic;
  signal bc_135 : std_logic;
  signal bc_136 : std_logic;
  signal bc_137 : std_logic;
  signal bc_138 : std_logic;
  signal bc_139 : std_logic;
  signal bc_140 : std_logic;
  signal bc_141 : std_logic;
  signal bc_142 : std_logic;
  signal bc_143 : std_logic;
  signal bc_144 : std_logic;
  signal bc_145 : std_logic;
  signal bc_146 : std_logic;
  signal bc_147 : std_logic;
  signal bc_148 : std_logic;
  signal bc_149 : std_logic;
  signal bc_150 : std_logic;
  signal bc_151 : std_logic;
  signal bc_152 : std_logic;
  signal bc_153 : std_logic;
  signal bc_154 : std_logic;
  signal bc_155 : std_logic;
  signal bc_156 : std_logic;
  signal bc_157 : std_logic;
  signal bc_158 : std_logic;
  signal bc_159 : std_logic;
  signal bc_160 : std_logic;
  signal bc_161 : std_logic;
  signal bc_162 : std_logic;
  signal bc_163 : std_logic;
  signal bc_164 : std_logic;
  signal bc_165 : std_logic;
  signal bc_166 : std_logic;
  signal bc_167 : std_logic;
  signal bc_168 : std_logic;
  signal bd_0 : std_logic;
  signal bd_1 : std_logic;
  signal bd_2 : std_logic;
  signal bd_3 : std_logic;
  signal bd_4 : std_logic;
  signal bd_5 : std_logic;
  signal bd_6 : std_logic;
  signal bd_7 : std_logic;
  signal bd_8 : std_logic;
  signal bd_9 : std_logic;
  signal bd_10 : std_logic;
  signal bd_11 : std_logic;
  signal bd_12 : std_logic;
  signal bd_13 : std_logic;
  signal bd_14 : std_logic;
  signal bd_15 : std_logic;
  signal bd_16 : std_logic;
  signal bd_17 : std_logic;
  signal bd_18 : std_logic;
  signal bd_19 : std_logic;
  signal bd_20 : std_logic;
  signal bd_21 : std_logic;
  signal bd_22 : std_logic;
  signal bd_23 : std_logic;
  signal bd_24 : std_logic;
  signal bd_25 : std_logic;
  signal bd_26 : std_logic;
  signal bd_27 : std_logic;
  signal bd_28 : std_logic;
  signal bd_29 : std_logic;
  signal bd_30 : std_logic;
  signal bd_31 : std_logic;
  signal bd_32 : std_logic;
  signal bd_33 : std_logic;
  signal bd_34 : std_logic;
  signal bd_35 : std_logic;
  signal bd_36 : std_logic;
  signal bd_37 : std_logic;
  signal bd_38 : std_logic;
  signal bd_39 : std_logic;
  signal bd_40 : std_logic;
  signal bd_41 : std_logic;
  signal bd_42 : std_logic;
  signal bd_43 : std_logic;
  signal bd_44 : std_logic;
  signal bd_45 : std_logic;
  signal bd_46 : std_logic;
  signal bd_47 : std_logic;
  signal bd_48 : std_logic;
  signal bd_49 : std_logic;
  signal bd_50 : std_logic;
  signal bd_51 : std_logic;
  signal bd_52 : std_logic;
  signal bd_53 : std_logic;
  signal bd_54 : std_logic;
  signal bd_55 : std_logic;
  signal bd_56 : std_logic;
  signal bd_57 : std_logic;
  signal bd_58 : std_logic;
  signal bd_59 : std_logic;
  signal bd_60 : std_logic;
  signal bd_61 : std_logic;
  signal bd_62 : std_logic;
  signal bd_63 : std_logic;
  signal bd_64 : std_logic;
  signal bd_65 : std_logic;
  signal bd_66 : std_logic;
  signal bd_67 : std_logic;
  signal bd_68 : std_logic;
  signal bd_69 : std_logic;
  signal bd_70 : std_logic;
  signal bd_71 : std_logic;
  signal bd_72 : std_logic;
  signal bd_73 : std_logic;
  signal bd_74 : std_logic;
  signal bd_75 : std_logic;
  signal bd_76 : std_logic;
  signal bd_77 : std_logic;
  signal bd_78 : std_logic;
  signal bd_79 : std_logic;
  signal bd_80 : std_logic;
  signal bd_81 : std_logic;
  signal bd_82 : std_logic;
  signal bd_83 : std_logic;
  signal bd_84 : std_logic;
  signal bd_85 : std_logic;
  signal bd_86 : std_logic;
  signal bd_87 : std_logic;
  signal bd_88 : std_logic;
  signal bd_89 : std_logic;
  signal bd_90 : std_logic;
  signal bd_91 : std_logic;
  signal bd_92 : std_logic;
  signal bd_93 : std_logic;
  signal bd_94 : std_logic;
  signal bd_95 : std_logic;
  signal bd_96 : std_logic;
  signal bd_97 : std_logic;
  signal bd_98 : std_logic;
  signal bd_99 : std_logic;
  signal bd_100 : std_logic;
  signal bd_101 : std_logic;
  signal bd_102 : std_logic;
  signal bd_103 : std_logic;
  signal bd_104 : std_logic;
  signal bd_105 : std_logic;
  signal bd_106 : std_logic;
  signal bd_107 : std_logic;
  signal bd_108 : std_logic;
  signal bd_109 : std_logic;
  signal bd_110 : std_logic;
  signal bd_111 : std_logic;
  signal bd_112 : std_logic;
  signal bd_113 : std_logic;
  signal bd_114 : std_logic;
  signal bd_115 : std_logic;
  signal bd_116 : std_logic;
  signal bd_117 : std_logic;
  signal bd_118 : std_logic;
  signal bd_119 : std_logic;
  signal bd_120 : std_logic;
  signal bd_121 : std_logic;
  signal bd_122 : std_logic;
  signal bd_123 : std_logic;
  signal bd_124 : std_logic;
  signal bd_125 : std_logic;
  signal bd_126 : std_logic;
  signal bd_127 : std_logic;
  signal bd_128 : std_logic;
  signal bd_129 : std_logic;
  signal bd_130 : std_logic;
  signal bd_131 : std_logic;
  signal bd_132 : std_logic;
  signal bd_133 : std_logic;
  signal bd_134 : std_logic;
  signal bd_135 : std_logic;
  signal bd_136 : std_logic;
  signal bd_137 : std_logic;
  signal bd_138 : std_logic;
  signal bd_139 : std_logic;
  signal bd_140 : std_logic;
  signal bd_141 : std_logic;
  signal bd_142 : std_logic;
  signal bd_143 : std_logic;
  signal bd_144 : std_logic;
  signal bd_145 : std_logic;
  signal bd_146 : std_logic;
  signal bd_147 : std_logic;
  signal bd_148 : std_logic;
  signal bd_149 : std_logic;
  signal bd_150 : std_logic;
  signal bd_151 : std_logic;
  signal bd_152 : std_logic;
  signal bd_153 : std_logic;
  signal bd_154 : std_logic;
  signal bd_155 : std_logic;
  signal bd_156 : std_logic;
  signal bd_157 : std_logic;
  signal bd_158 : std_logic;
  signal bd_159 : std_logic;
  signal bd_160 : std_logic;
  signal bd_161 : std_logic;
  signal bd_162 : std_logic;
  signal bd_163 : std_logic;
  signal bd_164 : std_logic;
  signal bd_165 : std_logic;
  signal bd_166 : std_logic;
  signal bd_167 : std_logic;
  signal bd_168 : std_logic;
begin
  dummy <= pkg_toStdLogic(false);
  a_0 <= pkg_extract(io_x_0,1);
  b_0 <= pkg_extract(io_x_0,0);
  c_0 <= pkg_extract(io_y_0,1);
  d_0 <= pkg_extract(io_y_0,0);
  a_1 <= pkg_extract(io_x_1,1);
  b_1 <= pkg_extract(io_x_1,0);
  c_1 <= pkg_extract(io_y_1,1);
  d_1 <= pkg_extract(io_y_1,0);
  a_2 <= pkg_extract(io_x_2,1);
  b_2 <= pkg_extract(io_x_2,0);
  c_2 <= pkg_extract(io_y_2,1);
  d_2 <= pkg_extract(io_y_2,0);
  a_3 <= pkg_extract(io_x_3,1);
  b_3 <= pkg_extract(io_x_3,0);
  c_3 <= pkg_extract(io_y_3,1);
  d_3 <= pkg_extract(io_y_3,0);
  a_4 <= pkg_extract(io_x_4,1);
  b_4 <= pkg_extract(io_x_4,0);
  c_4 <= pkg_extract(io_y_4,1);
  d_4 <= pkg_extract(io_y_4,0);
  a_5 <= pkg_extract(io_x_5,1);
  b_5 <= pkg_extract(io_x_5,0);
  c_5 <= pkg_extract(io_y_5,1);
  d_5 <= pkg_extract(io_y_5,0);
  a_6 <= pkg_extract(io_x_6,1);
  b_6 <= pkg_extract(io_x_6,0);
  c_6 <= pkg_extract(io_y_6,1);
  d_6 <= pkg_extract(io_y_6,0);
  a_7 <= pkg_extract(io_x_7,1);
  b_7 <= pkg_extract(io_x_7,0);
  c_7 <= pkg_extract(io_y_7,1);
  d_7 <= pkg_extract(io_y_7,0);
  a_8 <= pkg_extract(io_x_8,1);
  b_8 <= pkg_extract(io_x_8,0);
  c_8 <= pkg_extract(io_y_8,1);
  d_8 <= pkg_extract(io_y_8,0);
  a_9 <= pkg_extract(io_x_9,1);
  b_9 <= pkg_extract(io_x_9,0);
  c_9 <= pkg_extract(io_y_9,1);
  d_9 <= pkg_extract(io_y_9,0);
  a_10 <= pkg_extract(io_x_10,1);
  b_10 <= pkg_extract(io_x_10,0);
  c_10 <= pkg_extract(io_y_10,1);
  d_10 <= pkg_extract(io_y_10,0);
  a_11 <= pkg_extract(io_x_11,1);
  b_11 <= pkg_extract(io_x_11,0);
  c_11 <= pkg_extract(io_y_11,1);
  d_11 <= pkg_extract(io_y_11,0);
  a_12 <= pkg_extract(io_x_12,1);
  b_12 <= pkg_extract(io_x_12,0);
  c_12 <= pkg_extract(io_y_12,1);
  d_12 <= pkg_extract(io_y_12,0);
  ac_0 <= (a_0 and c_0);
  ad_0 <= (a_0 and d_0);
  bc_0 <= (b_0 and c_0);
  bd_0 <= (b_0 and d_0);
  ac_1 <= (a_0 and c_1);
  ad_1 <= (a_0 and d_1);
  bc_1 <= (b_0 and c_1);
  bd_1 <= (b_0 and d_1);
  ac_2 <= (a_0 and c_2);
  ad_2 <= (a_0 and d_2);
  bc_2 <= (b_0 and c_2);
  bd_2 <= (b_0 and d_2);
  ac_3 <= (a_0 and c_3);
  ad_3 <= (a_0 and d_3);
  bc_3 <= (b_0 and c_3);
  bd_3 <= (b_0 and d_3);
  ac_4 <= (a_0 and c_4);
  ad_4 <= (a_0 and d_4);
  bc_4 <= (b_0 and c_4);
  bd_4 <= (b_0 and d_4);
  ac_5 <= (a_0 and c_5);
  ad_5 <= (a_0 and d_5);
  bc_5 <= (b_0 and c_5);
  bd_5 <= (b_0 and d_5);
  ac_6 <= (a_0 and c_6);
  ad_6 <= (a_0 and d_6);
  bc_6 <= (b_0 and c_6);
  bd_6 <= (b_0 and d_6);
  ac_7 <= (a_0 and c_7);
  ad_7 <= (a_0 and d_7);
  bc_7 <= (b_0 and c_7);
  bd_7 <= (b_0 and d_7);
  ac_8 <= (a_0 and c_8);
  ad_8 <= (a_0 and d_8);
  bc_8 <= (b_0 and c_8);
  bd_8 <= (b_0 and d_8);
  ac_9 <= (a_0 and c_9);
  ad_9 <= (a_0 and d_9);
  bc_9 <= (b_0 and c_9);
  bd_9 <= (b_0 and d_9);
  ac_10 <= (a_0 and c_10);
  ad_10 <= (a_0 and d_10);
  bc_10 <= (b_0 and c_10);
  bd_10 <= (b_0 and d_10);
  ac_11 <= (a_0 and c_11);
  ad_11 <= (a_0 and d_11);
  bc_11 <= (b_0 and c_11);
  bd_11 <= (b_0 and d_11);
  ac_12 <= (a_0 and c_12);
  ad_12 <= (a_0 and d_12);
  bc_12 <= (b_0 and c_12);
  bd_12 <= (b_0 and d_12);
  ac_13 <= (a_1 and c_0);
  ad_13 <= (a_1 and d_0);
  bc_13 <= (b_1 and c_0);
  bd_13 <= (b_1 and d_0);
  ac_14 <= (a_1 and c_1);
  ad_14 <= (a_1 and d_1);
  bc_14 <= (b_1 and c_1);
  bd_14 <= (b_1 and d_1);
  ac_15 <= (a_1 and c_2);
  ad_15 <= (a_1 and d_2);
  bc_15 <= (b_1 and c_2);
  bd_15 <= (b_1 and d_2);
  ac_16 <= (a_1 and c_3);
  ad_16 <= (a_1 and d_3);
  bc_16 <= (b_1 and c_3);
  bd_16 <= (b_1 and d_3);
  ac_17 <= (a_1 and c_4);
  ad_17 <= (a_1 and d_4);
  bc_17 <= (b_1 and c_4);
  bd_17 <= (b_1 and d_4);
  ac_18 <= (a_1 and c_5);
  ad_18 <= (a_1 and d_5);
  bc_18 <= (b_1 and c_5);
  bd_18 <= (b_1 and d_5);
  ac_19 <= (a_1 and c_6);
  ad_19 <= (a_1 and d_6);
  bc_19 <= (b_1 and c_6);
  bd_19 <= (b_1 and d_6);
  ac_20 <= (a_1 and c_7);
  ad_20 <= (a_1 and d_7);
  bc_20 <= (b_1 and c_7);
  bd_20 <= (b_1 and d_7);
  ac_21 <= (a_1 and c_8);
  ad_21 <= (a_1 and d_8);
  bc_21 <= (b_1 and c_8);
  bd_21 <= (b_1 and d_8);
  ac_22 <= (a_1 and c_9);
  ad_22 <= (a_1 and d_9);
  bc_22 <= (b_1 and c_9);
  bd_22 <= (b_1 and d_9);
  ac_23 <= (a_1 and c_10);
  ad_23 <= (a_1 and d_10);
  bc_23 <= (b_1 and c_10);
  bd_23 <= (b_1 and d_10);
  ac_24 <= (a_1 and c_11);
  ad_24 <= (a_1 and d_11);
  bc_24 <= (b_1 and c_11);
  bd_24 <= (b_1 and d_11);
  ac_25 <= (a_1 and c_12);
  ad_25 <= (a_1 and d_12);
  bc_25 <= (b_1 and c_12);
  bd_25 <= (b_1 and d_12);
  ac_26 <= (a_2 and c_0);
  ad_26 <= (a_2 and d_0);
  bc_26 <= (b_2 and c_0);
  bd_26 <= (b_2 and d_0);
  ac_27 <= (a_2 and c_1);
  ad_27 <= (a_2 and d_1);
  bc_27 <= (b_2 and c_1);
  bd_27 <= (b_2 and d_1);
  ac_28 <= (a_2 and c_2);
  ad_28 <= (a_2 and d_2);
  bc_28 <= (b_2 and c_2);
  bd_28 <= (b_2 and d_2);
  ac_29 <= (a_2 and c_3);
  ad_29 <= (a_2 and d_3);
  bc_29 <= (b_2 and c_3);
  bd_29 <= (b_2 and d_3);
  ac_30 <= (a_2 and c_4);
  ad_30 <= (a_2 and d_4);
  bc_30 <= (b_2 and c_4);
  bd_30 <= (b_2 and d_4);
  ac_31 <= (a_2 and c_5);
  ad_31 <= (a_2 and d_5);
  bc_31 <= (b_2 and c_5);
  bd_31 <= (b_2 and d_5);
  ac_32 <= (a_2 and c_6);
  ad_32 <= (a_2 and d_6);
  bc_32 <= (b_2 and c_6);
  bd_32 <= (b_2 and d_6);
  ac_33 <= (a_2 and c_7);
  ad_33 <= (a_2 and d_7);
  bc_33 <= (b_2 and c_7);
  bd_33 <= (b_2 and d_7);
  ac_34 <= (a_2 and c_8);
  ad_34 <= (a_2 and d_8);
  bc_34 <= (b_2 and c_8);
  bd_34 <= (b_2 and d_8);
  ac_35 <= (a_2 and c_9);
  ad_35 <= (a_2 and d_9);
  bc_35 <= (b_2 and c_9);
  bd_35 <= (b_2 and d_9);
  ac_36 <= (a_2 and c_10);
  ad_36 <= (a_2 and d_10);
  bc_36 <= (b_2 and c_10);
  bd_36 <= (b_2 and d_10);
  ac_37 <= (a_2 and c_11);
  ad_37 <= (a_2 and d_11);
  bc_37 <= (b_2 and c_11);
  bd_37 <= (b_2 and d_11);
  ac_38 <= (a_2 and c_12);
  ad_38 <= (a_2 and d_12);
  bc_38 <= (b_2 and c_12);
  bd_38 <= (b_2 and d_12);
  ac_39 <= (a_3 and c_0);
  ad_39 <= (a_3 and d_0);
  bc_39 <= (b_3 and c_0);
  bd_39 <= (b_3 and d_0);
  ac_40 <= (a_3 and c_1);
  ad_40 <= (a_3 and d_1);
  bc_40 <= (b_3 and c_1);
  bd_40 <= (b_3 and d_1);
  ac_41 <= (a_3 and c_2);
  ad_41 <= (a_3 and d_2);
  bc_41 <= (b_3 and c_2);
  bd_41 <= (b_3 and d_2);
  ac_42 <= (a_3 and c_3);
  ad_42 <= (a_3 and d_3);
  bc_42 <= (b_3 and c_3);
  bd_42 <= (b_3 and d_3);
  ac_43 <= (a_3 and c_4);
  ad_43 <= (a_3 and d_4);
  bc_43 <= (b_3 and c_4);
  bd_43 <= (b_3 and d_4);
  ac_44 <= (a_3 and c_5);
  ad_44 <= (a_3 and d_5);
  bc_44 <= (b_3 and c_5);
  bd_44 <= (b_3 and d_5);
  ac_45 <= (a_3 and c_6);
  ad_45 <= (a_3 and d_6);
  bc_45 <= (b_3 and c_6);
  bd_45 <= (b_3 and d_6);
  ac_46 <= (a_3 and c_7);
  ad_46 <= (a_3 and d_7);
  bc_46 <= (b_3 and c_7);
  bd_46 <= (b_3 and d_7);
  ac_47 <= (a_3 and c_8);
  ad_47 <= (a_3 and d_8);
  bc_47 <= (b_3 and c_8);
  bd_47 <= (b_3 and d_8);
  ac_48 <= (a_3 and c_9);
  ad_48 <= (a_3 and d_9);
  bc_48 <= (b_3 and c_9);
  bd_48 <= (b_3 and d_9);
  ac_49 <= (a_3 and c_10);
  ad_49 <= (a_3 and d_10);
  bc_49 <= (b_3 and c_10);
  bd_49 <= (b_3 and d_10);
  ac_50 <= (a_3 and c_11);
  ad_50 <= (a_3 and d_11);
  bc_50 <= (b_3 and c_11);
  bd_50 <= (b_3 and d_11);
  ac_51 <= (a_3 and c_12);
  ad_51 <= (a_3 and d_12);
  bc_51 <= (b_3 and c_12);
  bd_51 <= (b_3 and d_12);
  ac_52 <= (a_4 and c_0);
  ad_52 <= (a_4 and d_0);
  bc_52 <= (b_4 and c_0);
  bd_52 <= (b_4 and d_0);
  ac_53 <= (a_4 and c_1);
  ad_53 <= (a_4 and d_1);
  bc_53 <= (b_4 and c_1);
  bd_53 <= (b_4 and d_1);
  ac_54 <= (a_4 and c_2);
  ad_54 <= (a_4 and d_2);
  bc_54 <= (b_4 and c_2);
  bd_54 <= (b_4 and d_2);
  ac_55 <= (a_4 and c_3);
  ad_55 <= (a_4 and d_3);
  bc_55 <= (b_4 and c_3);
  bd_55 <= (b_4 and d_3);
  ac_56 <= (a_4 and c_4);
  ad_56 <= (a_4 and d_4);
  bc_56 <= (b_4 and c_4);
  bd_56 <= (b_4 and d_4);
  ac_57 <= (a_4 and c_5);
  ad_57 <= (a_4 and d_5);
  bc_57 <= (b_4 and c_5);
  bd_57 <= (b_4 and d_5);
  ac_58 <= (a_4 and c_6);
  ad_58 <= (a_4 and d_6);
  bc_58 <= (b_4 and c_6);
  bd_58 <= (b_4 and d_6);
  ac_59 <= (a_4 and c_7);
  ad_59 <= (a_4 and d_7);
  bc_59 <= (b_4 and c_7);
  bd_59 <= (b_4 and d_7);
  ac_60 <= (a_4 and c_8);
  ad_60 <= (a_4 and d_8);
  bc_60 <= (b_4 and c_8);
  bd_60 <= (b_4 and d_8);
  ac_61 <= (a_4 and c_9);
  ad_61 <= (a_4 and d_9);
  bc_61 <= (b_4 and c_9);
  bd_61 <= (b_4 and d_9);
  ac_62 <= (a_4 and c_10);
  ad_62 <= (a_4 and d_10);
  bc_62 <= (b_4 and c_10);
  bd_62 <= (b_4 and d_10);
  ac_63 <= (a_4 and c_11);
  ad_63 <= (a_4 and d_11);
  bc_63 <= (b_4 and c_11);
  bd_63 <= (b_4 and d_11);
  ac_64 <= (a_4 and c_12);
  ad_64 <= (a_4 and d_12);
  bc_64 <= (b_4 and c_12);
  bd_64 <= (b_4 and d_12);
  ac_65 <= (a_5 and c_0);
  ad_65 <= (a_5 and d_0);
  bc_65 <= (b_5 and c_0);
  bd_65 <= (b_5 and d_0);
  ac_66 <= (a_5 and c_1);
  ad_66 <= (a_5 and d_1);
  bc_66 <= (b_5 and c_1);
  bd_66 <= (b_5 and d_1);
  ac_67 <= (a_5 and c_2);
  ad_67 <= (a_5 and d_2);
  bc_67 <= (b_5 and c_2);
  bd_67 <= (b_5 and d_2);
  ac_68 <= (a_5 and c_3);
  ad_68 <= (a_5 and d_3);
  bc_68 <= (b_5 and c_3);
  bd_68 <= (b_5 and d_3);
  ac_69 <= (a_5 and c_4);
  ad_69 <= (a_5 and d_4);
  bc_69 <= (b_5 and c_4);
  bd_69 <= (b_5 and d_4);
  ac_70 <= (a_5 and c_5);
  ad_70 <= (a_5 and d_5);
  bc_70 <= (b_5 and c_5);
  bd_70 <= (b_5 and d_5);
  ac_71 <= (a_5 and c_6);
  ad_71 <= (a_5 and d_6);
  bc_71 <= (b_5 and c_6);
  bd_71 <= (b_5 and d_6);
  ac_72 <= (a_5 and c_7);
  ad_72 <= (a_5 and d_7);
  bc_72 <= (b_5 and c_7);
  bd_72 <= (b_5 and d_7);
  ac_73 <= (a_5 and c_8);
  ad_73 <= (a_5 and d_8);
  bc_73 <= (b_5 and c_8);
  bd_73 <= (b_5 and d_8);
  ac_74 <= (a_5 and c_9);
  ad_74 <= (a_5 and d_9);
  bc_74 <= (b_5 and c_9);
  bd_74 <= (b_5 and d_9);
  ac_75 <= (a_5 and c_10);
  ad_75 <= (a_5 and d_10);
  bc_75 <= (b_5 and c_10);
  bd_75 <= (b_5 and d_10);
  ac_76 <= (a_5 and c_11);
  ad_76 <= (a_5 and d_11);
  bc_76 <= (b_5 and c_11);
  bd_76 <= (b_5 and d_11);
  ac_77 <= (a_5 and c_12);
  ad_77 <= (a_5 and d_12);
  bc_77 <= (b_5 and c_12);
  bd_77 <= (b_5 and d_12);
  ac_78 <= (a_6 and c_0);
  ad_78 <= (a_6 and d_0);
  bc_78 <= (b_6 and c_0);
  bd_78 <= (b_6 and d_0);
  ac_79 <= (a_6 and c_1);
  ad_79 <= (a_6 and d_1);
  bc_79 <= (b_6 and c_1);
  bd_79 <= (b_6 and d_1);
  ac_80 <= (a_6 and c_2);
  ad_80 <= (a_6 and d_2);
  bc_80 <= (b_6 and c_2);
  bd_80 <= (b_6 and d_2);
  ac_81 <= (a_6 and c_3);
  ad_81 <= (a_6 and d_3);
  bc_81 <= (b_6 and c_3);
  bd_81 <= (b_6 and d_3);
  ac_82 <= (a_6 and c_4);
  ad_82 <= (a_6 and d_4);
  bc_82 <= (b_6 and c_4);
  bd_82 <= (b_6 and d_4);
  ac_83 <= (a_6 and c_5);
  ad_83 <= (a_6 and d_5);
  bc_83 <= (b_6 and c_5);
  bd_83 <= (b_6 and d_5);
  ac_84 <= (a_6 and c_6);
  ad_84 <= (a_6 and d_6);
  bc_84 <= (b_6 and c_6);
  bd_84 <= (b_6 and d_6);
  ac_85 <= (a_6 and c_7);
  ad_85 <= (a_6 and d_7);
  bc_85 <= (b_6 and c_7);
  bd_85 <= (b_6 and d_7);
  ac_86 <= (a_6 and c_8);
  ad_86 <= (a_6 and d_8);
  bc_86 <= (b_6 and c_8);
  bd_86 <= (b_6 and d_8);
  ac_87 <= (a_6 and c_9);
  ad_87 <= (a_6 and d_9);
  bc_87 <= (b_6 and c_9);
  bd_87 <= (b_6 and d_9);
  ac_88 <= (a_6 and c_10);
  ad_88 <= (a_6 and d_10);
  bc_88 <= (b_6 and c_10);
  bd_88 <= (b_6 and d_10);
  ac_89 <= (a_6 and c_11);
  ad_89 <= (a_6 and d_11);
  bc_89 <= (b_6 and c_11);
  bd_89 <= (b_6 and d_11);
  ac_90 <= (a_6 and c_12);
  ad_90 <= (a_6 and d_12);
  bc_90 <= (b_6 and c_12);
  bd_90 <= (b_6 and d_12);
  ac_91 <= (a_7 and c_0);
  ad_91 <= (a_7 and d_0);
  bc_91 <= (b_7 and c_0);
  bd_91 <= (b_7 and d_0);
  ac_92 <= (a_7 and c_1);
  ad_92 <= (a_7 and d_1);
  bc_92 <= (b_7 and c_1);
  bd_92 <= (b_7 and d_1);
  ac_93 <= (a_7 and c_2);
  ad_93 <= (a_7 and d_2);
  bc_93 <= (b_7 and c_2);
  bd_93 <= (b_7 and d_2);
  ac_94 <= (a_7 and c_3);
  ad_94 <= (a_7 and d_3);
  bc_94 <= (b_7 and c_3);
  bd_94 <= (b_7 and d_3);
  ac_95 <= (a_7 and c_4);
  ad_95 <= (a_7 and d_4);
  bc_95 <= (b_7 and c_4);
  bd_95 <= (b_7 and d_4);
  ac_96 <= (a_7 and c_5);
  ad_96 <= (a_7 and d_5);
  bc_96 <= (b_7 and c_5);
  bd_96 <= (b_7 and d_5);
  ac_97 <= (a_7 and c_6);
  ad_97 <= (a_7 and d_6);
  bc_97 <= (b_7 and c_6);
  bd_97 <= (b_7 and d_6);
  ac_98 <= (a_7 and c_7);
  ad_98 <= (a_7 and d_7);
  bc_98 <= (b_7 and c_7);
  bd_98 <= (b_7 and d_7);
  ac_99 <= (a_7 and c_8);
  ad_99 <= (a_7 and d_8);
  bc_99 <= (b_7 and c_8);
  bd_99 <= (b_7 and d_8);
  ac_100 <= (a_7 and c_9);
  ad_100 <= (a_7 and d_9);
  bc_100 <= (b_7 and c_9);
  bd_100 <= (b_7 and d_9);
  ac_101 <= (a_7 and c_10);
  ad_101 <= (a_7 and d_10);
  bc_101 <= (b_7 and c_10);
  bd_101 <= (b_7 and d_10);
  ac_102 <= (a_7 and c_11);
  ad_102 <= (a_7 and d_11);
  bc_102 <= (b_7 and c_11);
  bd_102 <= (b_7 and d_11);
  ac_103 <= (a_7 and c_12);
  ad_103 <= (a_7 and d_12);
  bc_103 <= (b_7 and c_12);
  bd_103 <= (b_7 and d_12);
  ac_104 <= (a_8 and c_0);
  ad_104 <= (a_8 and d_0);
  bc_104 <= (b_8 and c_0);
  bd_104 <= (b_8 and d_0);
  ac_105 <= (a_8 and c_1);
  ad_105 <= (a_8 and d_1);
  bc_105 <= (b_8 and c_1);
  bd_105 <= (b_8 and d_1);
  ac_106 <= (a_8 and c_2);
  ad_106 <= (a_8 and d_2);
  bc_106 <= (b_8 and c_2);
  bd_106 <= (b_8 and d_2);
  ac_107 <= (a_8 and c_3);
  ad_107 <= (a_8 and d_3);
  bc_107 <= (b_8 and c_3);
  bd_107 <= (b_8 and d_3);
  ac_108 <= (a_8 and c_4);
  ad_108 <= (a_8 and d_4);
  bc_108 <= (b_8 and c_4);
  bd_108 <= (b_8 and d_4);
  ac_109 <= (a_8 and c_5);
  ad_109 <= (a_8 and d_5);
  bc_109 <= (b_8 and c_5);
  bd_109 <= (b_8 and d_5);
  ac_110 <= (a_8 and c_6);
  ad_110 <= (a_8 and d_6);
  bc_110 <= (b_8 and c_6);
  bd_110 <= (b_8 and d_6);
  ac_111 <= (a_8 and c_7);
  ad_111 <= (a_8 and d_7);
  bc_111 <= (b_8 and c_7);
  bd_111 <= (b_8 and d_7);
  ac_112 <= (a_8 and c_8);
  ad_112 <= (a_8 and d_8);
  bc_112 <= (b_8 and c_8);
  bd_112 <= (b_8 and d_8);
  ac_113 <= (a_8 and c_9);
  ad_113 <= (a_8 and d_9);
  bc_113 <= (b_8 and c_9);
  bd_113 <= (b_8 and d_9);
  ac_114 <= (a_8 and c_10);
  ad_114 <= (a_8 and d_10);
  bc_114 <= (b_8 and c_10);
  bd_114 <= (b_8 and d_10);
  ac_115 <= (a_8 and c_11);
  ad_115 <= (a_8 and d_11);
  bc_115 <= (b_8 and c_11);
  bd_115 <= (b_8 and d_11);
  ac_116 <= (a_8 and c_12);
  ad_116 <= (a_8 and d_12);
  bc_116 <= (b_8 and c_12);
  bd_116 <= (b_8 and d_12);
  ac_117 <= (a_9 and c_0);
  ad_117 <= (a_9 and d_0);
  bc_117 <= (b_9 and c_0);
  bd_117 <= (b_9 and d_0);
  ac_118 <= (a_9 and c_1);
  ad_118 <= (a_9 and d_1);
  bc_118 <= (b_9 and c_1);
  bd_118 <= (b_9 and d_1);
  ac_119 <= (a_9 and c_2);
  ad_119 <= (a_9 and d_2);
  bc_119 <= (b_9 and c_2);
  bd_119 <= (b_9 and d_2);
  ac_120 <= (a_9 and c_3);
  ad_120 <= (a_9 and d_3);
  bc_120 <= (b_9 and c_3);
  bd_120 <= (b_9 and d_3);
  ac_121 <= (a_9 and c_4);
  ad_121 <= (a_9 and d_4);
  bc_121 <= (b_9 and c_4);
  bd_121 <= (b_9 and d_4);
  ac_122 <= (a_9 and c_5);
  ad_122 <= (a_9 and d_5);
  bc_122 <= (b_9 and c_5);
  bd_122 <= (b_9 and d_5);
  ac_123 <= (a_9 and c_6);
  ad_123 <= (a_9 and d_6);
  bc_123 <= (b_9 and c_6);
  bd_123 <= (b_9 and d_6);
  ac_124 <= (a_9 and c_7);
  ad_124 <= (a_9 and d_7);
  bc_124 <= (b_9 and c_7);
  bd_124 <= (b_9 and d_7);
  ac_125 <= (a_9 and c_8);
  ad_125 <= (a_9 and d_8);
  bc_125 <= (b_9 and c_8);
  bd_125 <= (b_9 and d_8);
  ac_126 <= (a_9 and c_9);
  ad_126 <= (a_9 and d_9);
  bc_126 <= (b_9 and c_9);
  bd_126 <= (b_9 and d_9);
  ac_127 <= (a_9 and c_10);
  ad_127 <= (a_9 and d_10);
  bc_127 <= (b_9 and c_10);
  bd_127 <= (b_9 and d_10);
  ac_128 <= (a_9 and c_11);
  ad_128 <= (a_9 and d_11);
  bc_128 <= (b_9 and c_11);
  bd_128 <= (b_9 and d_11);
  ac_129 <= (a_9 and c_12);
  ad_129 <= (a_9 and d_12);
  bc_129 <= (b_9 and c_12);
  bd_129 <= (b_9 and d_12);
  ac_130 <= (a_10 and c_0);
  ad_130 <= (a_10 and d_0);
  bc_130 <= (b_10 and c_0);
  bd_130 <= (b_10 and d_0);
  ac_131 <= (a_10 and c_1);
  ad_131 <= (a_10 and d_1);
  bc_131 <= (b_10 and c_1);
  bd_131 <= (b_10 and d_1);
  ac_132 <= (a_10 and c_2);
  ad_132 <= (a_10 and d_2);
  bc_132 <= (b_10 and c_2);
  bd_132 <= (b_10 and d_2);
  ac_133 <= (a_10 and c_3);
  ad_133 <= (a_10 and d_3);
  bc_133 <= (b_10 and c_3);
  bd_133 <= (b_10 and d_3);
  ac_134 <= (a_10 and c_4);
  ad_134 <= (a_10 and d_4);
  bc_134 <= (b_10 and c_4);
  bd_134 <= (b_10 and d_4);
  ac_135 <= (a_10 and c_5);
  ad_135 <= (a_10 and d_5);
  bc_135 <= (b_10 and c_5);
  bd_135 <= (b_10 and d_5);
  ac_136 <= (a_10 and c_6);
  ad_136 <= (a_10 and d_6);
  bc_136 <= (b_10 and c_6);
  bd_136 <= (b_10 and d_6);
  ac_137 <= (a_10 and c_7);
  ad_137 <= (a_10 and d_7);
  bc_137 <= (b_10 and c_7);
  bd_137 <= (b_10 and d_7);
  ac_138 <= (a_10 and c_8);
  ad_138 <= (a_10 and d_8);
  bc_138 <= (b_10 and c_8);
  bd_138 <= (b_10 and d_8);
  ac_139 <= (a_10 and c_9);
  ad_139 <= (a_10 and d_9);
  bc_139 <= (b_10 and c_9);
  bd_139 <= (b_10 and d_9);
  ac_140 <= (a_10 and c_10);
  ad_140 <= (a_10 and d_10);
  bc_140 <= (b_10 and c_10);
  bd_140 <= (b_10 and d_10);
  ac_141 <= (a_10 and c_11);
  ad_141 <= (a_10 and d_11);
  bc_141 <= (b_10 and c_11);
  bd_141 <= (b_10 and d_11);
  ac_142 <= (a_10 and c_12);
  ad_142 <= (a_10 and d_12);
  bc_142 <= (b_10 and c_12);
  bd_142 <= (b_10 and d_12);
  ac_143 <= (a_11 and c_0);
  ad_143 <= (a_11 and d_0);
  bc_143 <= (b_11 and c_0);
  bd_143 <= (b_11 and d_0);
  ac_144 <= (a_11 and c_1);
  ad_144 <= (a_11 and d_1);
  bc_144 <= (b_11 and c_1);
  bd_144 <= (b_11 and d_1);
  ac_145 <= (a_11 and c_2);
  ad_145 <= (a_11 and d_2);
  bc_145 <= (b_11 and c_2);
  bd_145 <= (b_11 and d_2);
  ac_146 <= (a_11 and c_3);
  ad_146 <= (a_11 and d_3);
  bc_146 <= (b_11 and c_3);
  bd_146 <= (b_11 and d_3);
  ac_147 <= (a_11 and c_4);
  ad_147 <= (a_11 and d_4);
  bc_147 <= (b_11 and c_4);
  bd_147 <= (b_11 and d_4);
  ac_148 <= (a_11 and c_5);
  ad_148 <= (a_11 and d_5);
  bc_148 <= (b_11 and c_5);
  bd_148 <= (b_11 and d_5);
  ac_149 <= (a_11 and c_6);
  ad_149 <= (a_11 and d_6);
  bc_149 <= (b_11 and c_6);
  bd_149 <= (b_11 and d_6);
  ac_150 <= (a_11 and c_7);
  ad_150 <= (a_11 and d_7);
  bc_150 <= (b_11 and c_7);
  bd_150 <= (b_11 and d_7);
  ac_151 <= (a_11 and c_8);
  ad_151 <= (a_11 and d_8);
  bc_151 <= (b_11 and c_8);
  bd_151 <= (b_11 and d_8);
  ac_152 <= (a_11 and c_9);
  ad_152 <= (a_11 and d_9);
  bc_152 <= (b_11 and c_9);
  bd_152 <= (b_11 and d_9);
  ac_153 <= (a_11 and c_10);
  ad_153 <= (a_11 and d_10);
  bc_153 <= (b_11 and c_10);
  bd_153 <= (b_11 and d_10);
  ac_154 <= (a_11 and c_11);
  ad_154 <= (a_11 and d_11);
  bc_154 <= (b_11 and c_11);
  bd_154 <= (b_11 and d_11);
  ac_155 <= (a_11 and c_12);
  ad_155 <= (a_11 and d_12);
  bc_155 <= (b_11 and c_12);
  bd_155 <= (b_11 and d_12);
  ac_156 <= (a_12 and c_0);
  ad_156 <= (a_12 and d_0);
  bc_156 <= (b_12 and c_0);
  bd_156 <= (b_12 and d_0);
  ac_157 <= (a_12 and c_1);
  ad_157 <= (a_12 and d_1);
  bc_157 <= (b_12 and c_1);
  bd_157 <= (b_12 and d_1);
  ac_158 <= (a_12 and c_2);
  ad_158 <= (a_12 and d_2);
  bc_158 <= (b_12 and c_2);
  bd_158 <= (b_12 and d_2);
  ac_159 <= (a_12 and c_3);
  ad_159 <= (a_12 and d_3);
  bc_159 <= (b_12 and c_3);
  bd_159 <= (b_12 and d_3);
  ac_160 <= (a_12 and c_4);
  ad_160 <= (a_12 and d_4);
  bc_160 <= (b_12 and c_4);
  bd_160 <= (b_12 and d_4);
  ac_161 <= (a_12 and c_5);
  ad_161 <= (a_12 and d_5);
  bc_161 <= (b_12 and c_5);
  bd_161 <= (b_12 and d_5);
  ac_162 <= (a_12 and c_6);
  ad_162 <= (a_12 and d_6);
  bc_162 <= (b_12 and c_6);
  bd_162 <= (b_12 and d_6);
  ac_163 <= (a_12 and c_7);
  ad_163 <= (a_12 and d_7);
  bc_163 <= (b_12 and c_7);
  bd_163 <= (b_12 and d_7);
  ac_164 <= (a_12 and c_8);
  ad_164 <= (a_12 and d_8);
  bc_164 <= (b_12 and c_8);
  bd_164 <= (b_12 and d_8);
  ac_165 <= (a_12 and c_9);
  ad_165 <= (a_12 and d_9);
  bc_165 <= (b_12 and c_9);
  bd_165 <= (b_12 and d_9);
  ac_166 <= (a_12 and c_10);
  ad_166 <= (a_12 and d_10);
  bc_166 <= (b_12 and c_10);
  bd_166 <= (b_12 and d_10);
  ac_167 <= (a_12 and c_11);
  ad_167 <= (a_12 and d_11);
  bc_167 <= (b_12 and c_11);
  bd_167 <= (b_12 and d_11);
  ac_168 <= (a_12 and c_12);
  ad_168 <= (a_12 and d_12);
  bc_168 <= (b_12 and c_12);
  bd_168 <= (b_12 and d_12);
  process(bc_0,ad_0,bd_0,bc_14,ad_14,bd_14,bc_28,ad_28,bd_28,bc_42,ad_42,bd_42,bc_56,ad_56,bd_56,bc_70,ad_70,bd_70,bc_84,ad_84,bd_84,bc_98,ad_98,bd_98,bc_112,ad_112,bd_112,bc_126,ad_126,bd_126,bc_140,ad_140,bd_140,bc_154,ad_154,bd_154,bc_168,ad_168,bd_168)
  begin
    e_0(12) <= ((bc_0 xor ad_0) xor bd_0);
    e_0(0) <= ((bc_14 xor ad_14) xor bd_14);
    e_0(1) <= ((bc_28 xor ad_28) xor bd_28);
    e_0(2) <= ((bc_42 xor ad_42) xor bd_42);
    e_0(3) <= ((bc_56 xor ad_56) xor bd_56);
    e_0(4) <= ((bc_70 xor ad_70) xor bd_70);
    e_0(5) <= ((bc_84 xor ad_84) xor bd_84);
    e_0(6) <= ((bc_98 xor ad_98) xor bd_98);
    e_0(7) <= ((bc_112 xor ad_112) xor bd_112);
    e_0(8) <= ((bc_126 xor ad_126) xor bd_126);
    e_0(9) <= ((bc_140 xor ad_140) xor bd_140);
    e_0(10) <= ((bc_154 xor ad_154) xor bd_154);
    e_0(11) <= ((bc_168 xor ad_168) xor bd_168);
  end process;

  process(bc_0,ad_0,ac_0,bc_14,ad_14,ac_14,bc_28,ad_28,ac_28,bc_42,ad_42,ac_42,bc_56,ad_56,ac_56,bc_70,ad_70,ac_70,bc_84,ad_84,ac_84,bc_98,ad_98,ac_98,bc_112,ad_112,ac_112,bc_126,ad_126,ac_126,bc_140,ad_140,ac_140,bc_154,ad_154,ac_154,bc_168,ad_168,ac_168)
  begin
    f_0(12) <= ((bc_0 xor ad_0) xor ac_0);
    f_0(0) <= ((bc_14 xor ad_14) xor ac_14);
    f_0(1) <= ((bc_28 xor ad_28) xor ac_28);
    f_0(2) <= ((bc_42 xor ad_42) xor ac_42);
    f_0(3) <= ((bc_56 xor ad_56) xor ac_56);
    f_0(4) <= ((bc_70 xor ad_70) xor ac_70);
    f_0(5) <= ((bc_84 xor ad_84) xor ac_84);
    f_0(6) <= ((bc_98 xor ad_98) xor ac_98);
    f_0(7) <= ((bc_112 xor ad_112) xor ac_112);
    f_0(8) <= ((bc_126 xor ad_126) xor ac_126);
    f_0(9) <= ((bc_140 xor ad_140) xor ac_140);
    f_0(10) <= ((bc_154 xor ad_154) xor ac_154);
    f_0(11) <= ((bc_168 xor ad_168) xor ac_168);
  end process;

  process(e_0,bc_15,ad_15,bd_15,bc_2,ad_2,bd_2,bc_1,ad_1,bd_1,bc_4,ad_4,bd_4,bc_3,ad_3,bd_3,bc_6,ad_6,bd_6,bc_5,ad_5,bd_5,bc_8,ad_8,bd_8,bc_7,ad_7,bd_7,bc_10,ad_10,bd_10,bc_9,ad_9,bd_9,bc_12,ad_12,bd_12,bc_11,ad_11,bd_11)
  begin
    e_1(0) <= (((pkg_extract(e_0,0) xor bc_15) xor ad_15) xor bd_15);
    e_1(1) <= (((pkg_extract(e_0,1) xor bc_2) xor ad_2) xor bd_2);
    e_1(2) <= (((pkg_extract(e_0,2) xor bc_1) xor ad_1) xor bd_1);
    e_1(3) <= (((pkg_extract(e_0,3) xor bc_4) xor ad_4) xor bd_4);
    e_1(4) <= (((pkg_extract(e_0,4) xor bc_3) xor ad_3) xor bd_3);
    e_1(5) <= (((pkg_extract(e_0,5) xor bc_6) xor ad_6) xor bd_6);
    e_1(6) <= (((pkg_extract(e_0,6) xor bc_5) xor ad_5) xor bd_5);
    e_1(7) <= (((pkg_extract(e_0,7) xor bc_8) xor ad_8) xor bd_8);
    e_1(8) <= (((pkg_extract(e_0,8) xor bc_7) xor ad_7) xor bd_7);
    e_1(9) <= (((pkg_extract(e_0,9) xor bc_10) xor ad_10) xor bd_10);
    e_1(10) <= (((pkg_extract(e_0,10) xor bc_9) xor ad_9) xor bd_9);
    e_1(11) <= (((pkg_extract(e_0,11) xor bc_12) xor ad_12) xor bd_12);
    e_1(12) <= (((pkg_extract(e_0,12) xor bc_11) xor ad_11) xor bd_11);
  end process;

  process(f_0,bc_15,ad_15,ac_15,bc_2,ad_2,ac_2,bc_1,ad_1,ac_1,bc_4,ad_4,ac_4,bc_3,ad_3,ac_3,bc_6,ad_6,ac_6,bc_5,ad_5,ac_5,bc_8,ad_8,ac_8,bc_7,ad_7,ac_7,bc_10,ad_10,ac_10,bc_9,ad_9,ac_9,bc_12,ad_12,ac_12,bc_11,ad_11,ac_11)
  begin
    f_1(0) <= (((pkg_extract(f_0,0) xor bc_15) xor ad_15) xor ac_15);
    f_1(1) <= (((pkg_extract(f_0,1) xor bc_2) xor ad_2) xor ac_2);
    f_1(2) <= (((pkg_extract(f_0,2) xor bc_1) xor ad_1) xor ac_1);
    f_1(3) <= (((pkg_extract(f_0,3) xor bc_4) xor ad_4) xor ac_4);
    f_1(4) <= (((pkg_extract(f_0,4) xor bc_3) xor ad_3) xor ac_3);
    f_1(5) <= (((pkg_extract(f_0,5) xor bc_6) xor ad_6) xor ac_6);
    f_1(6) <= (((pkg_extract(f_0,6) xor bc_5) xor ad_5) xor ac_5);
    f_1(7) <= (((pkg_extract(f_0,7) xor bc_8) xor ad_8) xor ac_8);
    f_1(8) <= (((pkg_extract(f_0,8) xor bc_7) xor ad_7) xor ac_7);
    f_1(9) <= (((pkg_extract(f_0,9) xor bc_10) xor ad_10) xor ac_10);
    f_1(10) <= (((pkg_extract(f_0,10) xor bc_9) xor ad_9) xor ac_9);
    f_1(11) <= (((pkg_extract(f_0,11) xor bc_12) xor ad_12) xor ac_12);
    f_1(12) <= (((pkg_extract(f_0,12) xor bc_11) xor ad_11) xor ac_11);
  end process;

  process(e_1,bc_27,ad_27,bd_27,bc_26,ad_26,bd_26,bc_13,ad_13,bd_13,bc_17,ad_17,bd_17,bc_16,ad_16,bd_16,bc_19,ad_19,bd_19,bc_18,ad_18,bd_18,bc_21,ad_21,bd_21,bc_20,ad_20,bd_20,bc_23,ad_23,bd_23,bc_22,ad_22,bd_22,bc_25,ad_25,bd_25,bc_24,ad_24,bd_24)
  begin
    e_2(0) <= (((pkg_extract(e_1,0) xor bc_27) xor ad_27) xor bd_27);
    e_2(1) <= (((pkg_extract(e_1,1) xor bc_26) xor ad_26) xor bd_26);
    e_2(2) <= (((pkg_extract(e_1,2) xor bc_13) xor ad_13) xor bd_13);
    e_2(3) <= (((pkg_extract(e_1,3) xor bc_17) xor ad_17) xor bd_17);
    e_2(4) <= (((pkg_extract(e_1,4) xor bc_16) xor ad_16) xor bd_16);
    e_2(5) <= (((pkg_extract(e_1,5) xor bc_19) xor ad_19) xor bd_19);
    e_2(6) <= (((pkg_extract(e_1,6) xor bc_18) xor ad_18) xor bd_18);
    e_2(7) <= (((pkg_extract(e_1,7) xor bc_21) xor ad_21) xor bd_21);
    e_2(8) <= (((pkg_extract(e_1,8) xor bc_20) xor ad_20) xor bd_20);
    e_2(9) <= (((pkg_extract(e_1,9) xor bc_23) xor ad_23) xor bd_23);
    e_2(10) <= (((pkg_extract(e_1,10) xor bc_22) xor ad_22) xor bd_22);
    e_2(11) <= (((pkg_extract(e_1,11) xor bc_25) xor ad_25) xor bd_25);
    e_2(12) <= (((pkg_extract(e_1,12) xor bc_24) xor ad_24) xor bd_24);
  end process;

  process(f_1,bc_27,ad_27,ac_27,bc_26,ad_26,ac_26,bc_13,ad_13,ac_13,bc_17,ad_17,ac_17,bc_16,ad_16,ac_16,bc_19,ad_19,ac_19,bc_18,ad_18,ac_18,bc_21,ad_21,ac_21,bc_20,ad_20,ac_20,bc_23,ad_23,ac_23,bc_22,ad_22,ac_22,bc_25,ad_25,ac_25,bc_24,ad_24,ac_24)
  begin
    f_2(0) <= (((pkg_extract(f_1,0) xor bc_27) xor ad_27) xor ac_27);
    f_2(1) <= (((pkg_extract(f_1,1) xor bc_26) xor ad_26) xor ac_26);
    f_2(2) <= (((pkg_extract(f_1,2) xor bc_13) xor ad_13) xor ac_13);
    f_2(3) <= (((pkg_extract(f_1,3) xor bc_17) xor ad_17) xor ac_17);
    f_2(4) <= (((pkg_extract(f_1,4) xor bc_16) xor ad_16) xor ac_16);
    f_2(5) <= (((pkg_extract(f_1,5) xor bc_19) xor ad_19) xor ac_19);
    f_2(6) <= (((pkg_extract(f_1,6) xor bc_18) xor ad_18) xor ac_18);
    f_2(7) <= (((pkg_extract(f_1,7) xor bc_21) xor ad_21) xor ac_21);
    f_2(8) <= (((pkg_extract(f_1,8) xor bc_20) xor ad_20) xor ac_20);
    f_2(9) <= (((pkg_extract(f_1,9) xor bc_23) xor ad_23) xor ac_23);
    f_2(10) <= (((pkg_extract(f_1,10) xor bc_22) xor ad_22) xor ac_22);
    f_2(11) <= (((pkg_extract(f_1,11) xor bc_25) xor ad_25) xor ac_25);
    f_2(12) <= (((pkg_extract(f_1,12) xor bc_24) xor ad_24) xor ac_24);
  end process;

  process(e_2,bc_40,ad_40,bd_40,bc_39,ad_39,bd_39,bc_43,ad_43,bd_43,bc_30,ad_30,bd_30,bc_29,ad_29,bd_29,bc_32,ad_32,bd_32,bc_31,ad_31,bd_31,bc_34,ad_34,bd_34,bc_33,ad_33,bd_33,bc_36,ad_36,bd_36,bc_35,ad_35,bd_35,bc_38,ad_38,bd_38,bc_37,ad_37,bd_37)
  begin
    e_3(0) <= (((pkg_extract(e_2,0) xor bc_40) xor ad_40) xor bd_40);
    e_3(1) <= (((pkg_extract(e_2,1) xor bc_39) xor ad_39) xor bd_39);
    e_3(2) <= (((pkg_extract(e_2,2) xor bc_43) xor ad_43) xor bd_43);
    e_3(3) <= (((pkg_extract(e_2,3) xor bc_30) xor ad_30) xor bd_30);
    e_3(4) <= (((pkg_extract(e_2,4) xor bc_29) xor ad_29) xor bd_29);
    e_3(5) <= (((pkg_extract(e_2,5) xor bc_32) xor ad_32) xor bd_32);
    e_3(6) <= (((pkg_extract(e_2,6) xor bc_31) xor ad_31) xor bd_31);
    e_3(7) <= (((pkg_extract(e_2,7) xor bc_34) xor ad_34) xor bd_34);
    e_3(8) <= (((pkg_extract(e_2,8) xor bc_33) xor ad_33) xor bd_33);
    e_3(9) <= (((pkg_extract(e_2,9) xor bc_36) xor ad_36) xor bd_36);
    e_3(10) <= (((pkg_extract(e_2,10) xor bc_35) xor ad_35) xor bd_35);
    e_3(11) <= (((pkg_extract(e_2,11) xor bc_38) xor ad_38) xor bd_38);
    e_3(12) <= (((pkg_extract(e_2,12) xor bc_37) xor ad_37) xor bd_37);
  end process;

  process(f_2,bc_40,ad_40,ac_40,bc_39,ad_39,ac_39,bc_43,ad_43,ac_43,bc_30,ad_30,ac_30,bc_29,ad_29,ac_29,bc_32,ad_32,ac_32,bc_31,ad_31,ac_31,bc_34,ad_34,ac_34,bc_33,ad_33,ac_33,bc_36,ad_36,ac_36,bc_35,ad_35,ac_35,bc_38,ad_38,ac_38,bc_37,ad_37,ac_37)
  begin
    f_3(0) <= (((pkg_extract(f_2,0) xor bc_40) xor ad_40) xor ac_40);
    f_3(1) <= (((pkg_extract(f_2,1) xor bc_39) xor ad_39) xor ac_39);
    f_3(2) <= (((pkg_extract(f_2,2) xor bc_43) xor ad_43) xor ac_43);
    f_3(3) <= (((pkg_extract(f_2,3) xor bc_30) xor ad_30) xor ac_30);
    f_3(4) <= (((pkg_extract(f_2,4) xor bc_29) xor ad_29) xor ac_29);
    f_3(5) <= (((pkg_extract(f_2,5) xor bc_32) xor ad_32) xor ac_32);
    f_3(6) <= (((pkg_extract(f_2,6) xor bc_31) xor ad_31) xor ac_31);
    f_3(7) <= (((pkg_extract(f_2,7) xor bc_34) xor ad_34) xor ac_34);
    f_3(8) <= (((pkg_extract(f_2,8) xor bc_33) xor ad_33) xor ac_33);
    f_3(9) <= (((pkg_extract(f_2,9) xor bc_36) xor ad_36) xor ac_36);
    f_3(10) <= (((pkg_extract(f_2,10) xor bc_35) xor ad_35) xor ac_35);
    f_3(11) <= (((pkg_extract(f_2,11) xor bc_38) xor ad_38) xor ac_38);
    f_3(12) <= (((pkg_extract(f_2,12) xor bc_37) xor ad_37) xor ac_37);
  end process;

  process(e_3,bc_53,ad_53,bd_53,bc_52,ad_52,bd_52,bc_55,ad_55,bd_55,bc_54,ad_54,bd_54,bc_41,ad_41,bd_41,bc_45,ad_45,bd_45,bc_44,ad_44,bd_44,bc_47,ad_47,bd_47,bc_46,ad_46,bd_46,bc_49,ad_49,bd_49,bc_48,ad_48,bd_48,bc_51,ad_51,bd_51,bc_50,ad_50,bd_50)
  begin
    e_4(0) <= (((pkg_extract(e_3,0) xor bc_53) xor ad_53) xor bd_53);
    e_4(1) <= (((pkg_extract(e_3,1) xor bc_52) xor ad_52) xor bd_52);
    e_4(2) <= (((pkg_extract(e_3,2) xor bc_55) xor ad_55) xor bd_55);
    e_4(3) <= (((pkg_extract(e_3,3) xor bc_54) xor ad_54) xor bd_54);
    e_4(4) <= (((pkg_extract(e_3,4) xor bc_41) xor ad_41) xor bd_41);
    e_4(5) <= (((pkg_extract(e_3,5) xor bc_45) xor ad_45) xor bd_45);
    e_4(6) <= (((pkg_extract(e_3,6) xor bc_44) xor ad_44) xor bd_44);
    e_4(7) <= (((pkg_extract(e_3,7) xor bc_47) xor ad_47) xor bd_47);
    e_4(8) <= (((pkg_extract(e_3,8) xor bc_46) xor ad_46) xor bd_46);
    e_4(9) <= (((pkg_extract(e_3,9) xor bc_49) xor ad_49) xor bd_49);
    e_4(10) <= (((pkg_extract(e_3,10) xor bc_48) xor ad_48) xor bd_48);
    e_4(11) <= (((pkg_extract(e_3,11) xor bc_51) xor ad_51) xor bd_51);
    e_4(12) <= (((pkg_extract(e_3,12) xor bc_50) xor ad_50) xor bd_50);
  end process;

  process(f_3,bc_53,ad_53,ac_53,bc_52,ad_52,ac_52,bc_55,ad_55,ac_55,bc_54,ad_54,ac_54,bc_41,ad_41,ac_41,bc_45,ad_45,ac_45,bc_44,ad_44,ac_44,bc_47,ad_47,ac_47,bc_46,ad_46,ac_46,bc_49,ad_49,ac_49,bc_48,ad_48,ac_48,bc_51,ad_51,ac_51,bc_50,ad_50,ac_50)
  begin
    f_4(0) <= (((pkg_extract(f_3,0) xor bc_53) xor ad_53) xor ac_53);
    f_4(1) <= (((pkg_extract(f_3,1) xor bc_52) xor ad_52) xor ac_52);
    f_4(2) <= (((pkg_extract(f_3,2) xor bc_55) xor ad_55) xor ac_55);
    f_4(3) <= (((pkg_extract(f_3,3) xor bc_54) xor ad_54) xor ac_54);
    f_4(4) <= (((pkg_extract(f_3,4) xor bc_41) xor ad_41) xor ac_41);
    f_4(5) <= (((pkg_extract(f_3,5) xor bc_45) xor ad_45) xor ac_45);
    f_4(6) <= (((pkg_extract(f_3,6) xor bc_44) xor ad_44) xor ac_44);
    f_4(7) <= (((pkg_extract(f_3,7) xor bc_47) xor ad_47) xor ac_47);
    f_4(8) <= (((pkg_extract(f_3,8) xor bc_46) xor ad_46) xor ac_46);
    f_4(9) <= (((pkg_extract(f_3,9) xor bc_49) xor ad_49) xor ac_49);
    f_4(10) <= (((pkg_extract(f_3,10) xor bc_48) xor ad_48) xor ac_48);
    f_4(11) <= (((pkg_extract(f_3,11) xor bc_51) xor ad_51) xor ac_51);
    f_4(12) <= (((pkg_extract(f_3,12) xor bc_50) xor ad_50) xor ac_50);
  end process;

  process(e_4,bc_66,ad_66,bd_66,bc_65,ad_65,bd_65,bc_68,ad_68,bd_68,bc_67,ad_67,bd_67,bc_71,ad_71,bd_71,bc_58,ad_58,bd_58,bc_57,ad_57,bd_57,bc_60,ad_60,bd_60,bc_59,ad_59,bd_59,bc_62,ad_62,bd_62,bc_61,ad_61,bd_61,bc_64,ad_64,bd_64,bc_63,ad_63,bd_63)
  begin
    e_5(0) <= (((pkg_extract(e_4,0) xor bc_66) xor ad_66) xor bd_66);
    e_5(1) <= (((pkg_extract(e_4,1) xor bc_65) xor ad_65) xor bd_65);
    e_5(2) <= (((pkg_extract(e_4,2) xor bc_68) xor ad_68) xor bd_68);
    e_5(3) <= (((pkg_extract(e_4,3) xor bc_67) xor ad_67) xor bd_67);
    e_5(4) <= (((pkg_extract(e_4,4) xor bc_71) xor ad_71) xor bd_71);
    e_5(5) <= (((pkg_extract(e_4,5) xor bc_58) xor ad_58) xor bd_58);
    e_5(6) <= (((pkg_extract(e_4,6) xor bc_57) xor ad_57) xor bd_57);
    e_5(7) <= (((pkg_extract(e_4,7) xor bc_60) xor ad_60) xor bd_60);
    e_5(8) <= (((pkg_extract(e_4,8) xor bc_59) xor ad_59) xor bd_59);
    e_5(9) <= (((pkg_extract(e_4,9) xor bc_62) xor ad_62) xor bd_62);
    e_5(10) <= (((pkg_extract(e_4,10) xor bc_61) xor ad_61) xor bd_61);
    e_5(11) <= (((pkg_extract(e_4,11) xor bc_64) xor ad_64) xor bd_64);
    e_5(12) <= (((pkg_extract(e_4,12) xor bc_63) xor ad_63) xor bd_63);
  end process;

  process(f_4,bc_66,ad_66,ac_66,bc_65,ad_65,ac_65,bc_68,ad_68,ac_68,bc_67,ad_67,ac_67,bc_71,ad_71,ac_71,bc_58,ad_58,ac_58,bc_57,ad_57,ac_57,bc_60,ad_60,ac_60,bc_59,ad_59,ac_59,bc_62,ad_62,ac_62,bc_61,ad_61,ac_61,bc_64,ad_64,ac_64,bc_63,ad_63,ac_63)
  begin
    f_5(0) <= (((pkg_extract(f_4,0) xor bc_66) xor ad_66) xor ac_66);
    f_5(1) <= (((pkg_extract(f_4,1) xor bc_65) xor ad_65) xor ac_65);
    f_5(2) <= (((pkg_extract(f_4,2) xor bc_68) xor ad_68) xor ac_68);
    f_5(3) <= (((pkg_extract(f_4,3) xor bc_67) xor ad_67) xor ac_67);
    f_5(4) <= (((pkg_extract(f_4,4) xor bc_71) xor ad_71) xor ac_71);
    f_5(5) <= (((pkg_extract(f_4,5) xor bc_58) xor ad_58) xor ac_58);
    f_5(6) <= (((pkg_extract(f_4,6) xor bc_57) xor ad_57) xor ac_57);
    f_5(7) <= (((pkg_extract(f_4,7) xor bc_60) xor ad_60) xor ac_60);
    f_5(8) <= (((pkg_extract(f_4,8) xor bc_59) xor ad_59) xor ac_59);
    f_5(9) <= (((pkg_extract(f_4,9) xor bc_62) xor ad_62) xor ac_62);
    f_5(10) <= (((pkg_extract(f_4,10) xor bc_61) xor ad_61) xor ac_61);
    f_5(11) <= (((pkg_extract(f_4,11) xor bc_64) xor ad_64) xor ac_64);
    f_5(12) <= (((pkg_extract(f_4,12) xor bc_63) xor ad_63) xor ac_63);
  end process;

  process(e_5,bc_79,ad_79,bd_79,bc_78,ad_78,bd_78,bc_81,ad_81,bd_81,bc_80,ad_80,bd_80,bc_83,ad_83,bd_83,bc_82,ad_82,bd_82,bc_69,ad_69,bd_69,bc_73,ad_73,bd_73,bc_72,ad_72,bd_72,bc_75,ad_75,bd_75,bc_74,ad_74,bd_74,bc_77,ad_77,bd_77,bc_76,ad_76,bd_76)
  begin
    e_6(0) <= (((pkg_extract(e_5,0) xor bc_79) xor ad_79) xor bd_79);
    e_6(1) <= (((pkg_extract(e_5,1) xor bc_78) xor ad_78) xor bd_78);
    e_6(2) <= (((pkg_extract(e_5,2) xor bc_81) xor ad_81) xor bd_81);
    e_6(3) <= (((pkg_extract(e_5,3) xor bc_80) xor ad_80) xor bd_80);
    e_6(4) <= (((pkg_extract(e_5,4) xor bc_83) xor ad_83) xor bd_83);
    e_6(5) <= (((pkg_extract(e_5,5) xor bc_82) xor ad_82) xor bd_82);
    e_6(6) <= (((pkg_extract(e_5,6) xor bc_69) xor ad_69) xor bd_69);
    e_6(7) <= (((pkg_extract(e_5,7) xor bc_73) xor ad_73) xor bd_73);
    e_6(8) <= (((pkg_extract(e_5,8) xor bc_72) xor ad_72) xor bd_72);
    e_6(9) <= (((pkg_extract(e_5,9) xor bc_75) xor ad_75) xor bd_75);
    e_6(10) <= (((pkg_extract(e_5,10) xor bc_74) xor ad_74) xor bd_74);
    e_6(11) <= (((pkg_extract(e_5,11) xor bc_77) xor ad_77) xor bd_77);
    e_6(12) <= (((pkg_extract(e_5,12) xor bc_76) xor ad_76) xor bd_76);
  end process;

  process(f_5,bc_79,ad_79,ac_79,bc_78,ad_78,ac_78,bc_81,ad_81,ac_81,bc_80,ad_80,ac_80,bc_83,ad_83,ac_83,bc_82,ad_82,ac_82,bc_69,ad_69,ac_69,bc_73,ad_73,ac_73,bc_72,ad_72,ac_72,bc_75,ad_75,ac_75,bc_74,ad_74,ac_74,bc_77,ad_77,ac_77,bc_76,ad_76,ac_76)
  begin
    f_6(0) <= (((pkg_extract(f_5,0) xor bc_79) xor ad_79) xor ac_79);
    f_6(1) <= (((pkg_extract(f_5,1) xor bc_78) xor ad_78) xor ac_78);
    f_6(2) <= (((pkg_extract(f_5,2) xor bc_81) xor ad_81) xor ac_81);
    f_6(3) <= (((pkg_extract(f_5,3) xor bc_80) xor ad_80) xor ac_80);
    f_6(4) <= (((pkg_extract(f_5,4) xor bc_83) xor ad_83) xor ac_83);
    f_6(5) <= (((pkg_extract(f_5,5) xor bc_82) xor ad_82) xor ac_82);
    f_6(6) <= (((pkg_extract(f_5,6) xor bc_69) xor ad_69) xor ac_69);
    f_6(7) <= (((pkg_extract(f_5,7) xor bc_73) xor ad_73) xor ac_73);
    f_6(8) <= (((pkg_extract(f_5,8) xor bc_72) xor ad_72) xor ac_72);
    f_6(9) <= (((pkg_extract(f_5,9) xor bc_75) xor ad_75) xor ac_75);
    f_6(10) <= (((pkg_extract(f_5,10) xor bc_74) xor ad_74) xor ac_74);
    f_6(11) <= (((pkg_extract(f_5,11) xor bc_77) xor ad_77) xor ac_77);
    f_6(12) <= (((pkg_extract(f_5,12) xor bc_76) xor ad_76) xor ac_76);
  end process;

  process(e_6,bc_92,ad_92,bd_92,bc_91,ad_91,bd_91,bc_94,ad_94,bd_94,bc_93,ad_93,bd_93,bc_96,ad_96,bd_96,bc_95,ad_95,bd_95,bc_99,ad_99,bd_99,bc_86,ad_86,bd_86,bc_85,ad_85,bd_85,bc_88,ad_88,bd_88,bc_87,ad_87,bd_87,bc_90,ad_90,bd_90,bc_89,ad_89,bd_89)
  begin
    e_7(0) <= (((pkg_extract(e_6,0) xor bc_92) xor ad_92) xor bd_92);
    e_7(1) <= (((pkg_extract(e_6,1) xor bc_91) xor ad_91) xor bd_91);
    e_7(2) <= (((pkg_extract(e_6,2) xor bc_94) xor ad_94) xor bd_94);
    e_7(3) <= (((pkg_extract(e_6,3) xor bc_93) xor ad_93) xor bd_93);
    e_7(4) <= (((pkg_extract(e_6,4) xor bc_96) xor ad_96) xor bd_96);
    e_7(5) <= (((pkg_extract(e_6,5) xor bc_95) xor ad_95) xor bd_95);
    e_7(6) <= (((pkg_extract(e_6,6) xor bc_99) xor ad_99) xor bd_99);
    e_7(7) <= (((pkg_extract(e_6,7) xor bc_86) xor ad_86) xor bd_86);
    e_7(8) <= (((pkg_extract(e_6,8) xor bc_85) xor ad_85) xor bd_85);
    e_7(9) <= (((pkg_extract(e_6,9) xor bc_88) xor ad_88) xor bd_88);
    e_7(10) <= (((pkg_extract(e_6,10) xor bc_87) xor ad_87) xor bd_87);
    e_7(11) <= (((pkg_extract(e_6,11) xor bc_90) xor ad_90) xor bd_90);
    e_7(12) <= (((pkg_extract(e_6,12) xor bc_89) xor ad_89) xor bd_89);
  end process;

  process(f_6,bc_92,ad_92,ac_92,bc_91,ad_91,ac_91,bc_94,ad_94,ac_94,bc_93,ad_93,ac_93,bc_96,ad_96,ac_96,bc_95,ad_95,ac_95,bc_99,ad_99,ac_99,bc_86,ad_86,ac_86,bc_85,ad_85,ac_85,bc_88,ad_88,ac_88,bc_87,ad_87,ac_87,bc_90,ad_90,ac_90,bc_89,ad_89,ac_89)
  begin
    f_7(0) <= (((pkg_extract(f_6,0) xor bc_92) xor ad_92) xor ac_92);
    f_7(1) <= (((pkg_extract(f_6,1) xor bc_91) xor ad_91) xor ac_91);
    f_7(2) <= (((pkg_extract(f_6,2) xor bc_94) xor ad_94) xor ac_94);
    f_7(3) <= (((pkg_extract(f_6,3) xor bc_93) xor ad_93) xor ac_93);
    f_7(4) <= (((pkg_extract(f_6,4) xor bc_96) xor ad_96) xor ac_96);
    f_7(5) <= (((pkg_extract(f_6,5) xor bc_95) xor ad_95) xor ac_95);
    f_7(6) <= (((pkg_extract(f_6,6) xor bc_99) xor ad_99) xor ac_99);
    f_7(7) <= (((pkg_extract(f_6,7) xor bc_86) xor ad_86) xor ac_86);
    f_7(8) <= (((pkg_extract(f_6,8) xor bc_85) xor ad_85) xor ac_85);
    f_7(9) <= (((pkg_extract(f_6,9) xor bc_88) xor ad_88) xor ac_88);
    f_7(10) <= (((pkg_extract(f_6,10) xor bc_87) xor ad_87) xor ac_87);
    f_7(11) <= (((pkg_extract(f_6,11) xor bc_90) xor ad_90) xor ac_90);
    f_7(12) <= (((pkg_extract(f_6,12) xor bc_89) xor ad_89) xor ac_89);
  end process;

  process(e_7,bc_105,ad_105,bd_105,bc_104,ad_104,bd_104,bc_107,ad_107,bd_107,bc_106,ad_106,bd_106,bc_109,ad_109,bd_109,bc_108,ad_108,bd_108,bc_111,ad_111,bd_111,bc_110,ad_110,bd_110,bc_97,ad_97,bd_97,bc_101,ad_101,bd_101,bc_100,ad_100,bd_100,bc_103,ad_103,bd_103,bc_102,ad_102,bd_102)
  begin
    e_8(0) <= (((pkg_extract(e_7,0) xor bc_105) xor ad_105) xor bd_105);
    e_8(1) <= (((pkg_extract(e_7,1) xor bc_104) xor ad_104) xor bd_104);
    e_8(2) <= (((pkg_extract(e_7,2) xor bc_107) xor ad_107) xor bd_107);
    e_8(3) <= (((pkg_extract(e_7,3) xor bc_106) xor ad_106) xor bd_106);
    e_8(4) <= (((pkg_extract(e_7,4) xor bc_109) xor ad_109) xor bd_109);
    e_8(5) <= (((pkg_extract(e_7,5) xor bc_108) xor ad_108) xor bd_108);
    e_8(6) <= (((pkg_extract(e_7,6) xor bc_111) xor ad_111) xor bd_111);
    e_8(7) <= (((pkg_extract(e_7,7) xor bc_110) xor ad_110) xor bd_110);
    e_8(8) <= (((pkg_extract(e_7,8) xor bc_97) xor ad_97) xor bd_97);
    e_8(9) <= (((pkg_extract(e_7,9) xor bc_101) xor ad_101) xor bd_101);
    e_8(10) <= (((pkg_extract(e_7,10) xor bc_100) xor ad_100) xor bd_100);
    e_8(11) <= (((pkg_extract(e_7,11) xor bc_103) xor ad_103) xor bd_103);
    e_8(12) <= (((pkg_extract(e_7,12) xor bc_102) xor ad_102) xor bd_102);
  end process;

  process(f_7,bc_105,ad_105,ac_105,bc_104,ad_104,ac_104,bc_107,ad_107,ac_107,bc_106,ad_106,ac_106,bc_109,ad_109,ac_109,bc_108,ad_108,ac_108,bc_111,ad_111,ac_111,bc_110,ad_110,ac_110,bc_97,ad_97,ac_97,bc_101,ad_101,ac_101,bc_100,ad_100,ac_100,bc_103,ad_103,ac_103,bc_102,ad_102,ac_102)
  begin
    f_8(0) <= (((pkg_extract(f_7,0) xor bc_105) xor ad_105) xor ac_105);
    f_8(1) <= (((pkg_extract(f_7,1) xor bc_104) xor ad_104) xor ac_104);
    f_8(2) <= (((pkg_extract(f_7,2) xor bc_107) xor ad_107) xor ac_107);
    f_8(3) <= (((pkg_extract(f_7,3) xor bc_106) xor ad_106) xor ac_106);
    f_8(4) <= (((pkg_extract(f_7,4) xor bc_109) xor ad_109) xor ac_109);
    f_8(5) <= (((pkg_extract(f_7,5) xor bc_108) xor ad_108) xor ac_108);
    f_8(6) <= (((pkg_extract(f_7,6) xor bc_111) xor ad_111) xor ac_111);
    f_8(7) <= (((pkg_extract(f_7,7) xor bc_110) xor ad_110) xor ac_110);
    f_8(8) <= (((pkg_extract(f_7,8) xor bc_97) xor ad_97) xor ac_97);
    f_8(9) <= (((pkg_extract(f_7,9) xor bc_101) xor ad_101) xor ac_101);
    f_8(10) <= (((pkg_extract(f_7,10) xor bc_100) xor ad_100) xor ac_100);
    f_8(11) <= (((pkg_extract(f_7,11) xor bc_103) xor ad_103) xor ac_103);
    f_8(12) <= (((pkg_extract(f_7,12) xor bc_102) xor ad_102) xor ac_102);
  end process;

  process(e_8,bc_118,ad_118,bd_118,bc_117,ad_117,bd_117,bc_120,ad_120,bd_120,bc_119,ad_119,bd_119,bc_122,ad_122,bd_122,bc_121,ad_121,bd_121,bc_124,ad_124,bd_124,bc_123,ad_123,bd_123,bc_127,ad_127,bd_127,bc_114,ad_114,bd_114,bc_113,ad_113,bd_113,bc_116,ad_116,bd_116,bc_115,ad_115,bd_115)
  begin
    e_9(0) <= (((pkg_extract(e_8,0) xor bc_118) xor ad_118) xor bd_118);
    e_9(1) <= (((pkg_extract(e_8,1) xor bc_117) xor ad_117) xor bd_117);
    e_9(2) <= (((pkg_extract(e_8,2) xor bc_120) xor ad_120) xor bd_120);
    e_9(3) <= (((pkg_extract(e_8,3) xor bc_119) xor ad_119) xor bd_119);
    e_9(4) <= (((pkg_extract(e_8,4) xor bc_122) xor ad_122) xor bd_122);
    e_9(5) <= (((pkg_extract(e_8,5) xor bc_121) xor ad_121) xor bd_121);
    e_9(6) <= (((pkg_extract(e_8,6) xor bc_124) xor ad_124) xor bd_124);
    e_9(7) <= (((pkg_extract(e_8,7) xor bc_123) xor ad_123) xor bd_123);
    e_9(8) <= (((pkg_extract(e_8,8) xor bc_127) xor ad_127) xor bd_127);
    e_9(9) <= (((pkg_extract(e_8,9) xor bc_114) xor ad_114) xor bd_114);
    e_9(10) <= (((pkg_extract(e_8,10) xor bc_113) xor ad_113) xor bd_113);
    e_9(11) <= (((pkg_extract(e_8,11) xor bc_116) xor ad_116) xor bd_116);
    e_9(12) <= (((pkg_extract(e_8,12) xor bc_115) xor ad_115) xor bd_115);
  end process;

  process(f_8,bc_118,ad_118,ac_118,bc_117,ad_117,ac_117,bc_120,ad_120,ac_120,bc_119,ad_119,ac_119,bc_122,ad_122,ac_122,bc_121,ad_121,ac_121,bc_124,ad_124,ac_124,bc_123,ad_123,ac_123,bc_127,ad_127,ac_127,bc_114,ad_114,ac_114,bc_113,ad_113,ac_113,bc_116,ad_116,ac_116,bc_115,ad_115,ac_115)
  begin
    f_9(0) <= (((pkg_extract(f_8,0) xor bc_118) xor ad_118) xor ac_118);
    f_9(1) <= (((pkg_extract(f_8,1) xor bc_117) xor ad_117) xor ac_117);
    f_9(2) <= (((pkg_extract(f_8,2) xor bc_120) xor ad_120) xor ac_120);
    f_9(3) <= (((pkg_extract(f_8,3) xor bc_119) xor ad_119) xor ac_119);
    f_9(4) <= (((pkg_extract(f_8,4) xor bc_122) xor ad_122) xor ac_122);
    f_9(5) <= (((pkg_extract(f_8,5) xor bc_121) xor ad_121) xor ac_121);
    f_9(6) <= (((pkg_extract(f_8,6) xor bc_124) xor ad_124) xor ac_124);
    f_9(7) <= (((pkg_extract(f_8,7) xor bc_123) xor ad_123) xor ac_123);
    f_9(8) <= (((pkg_extract(f_8,8) xor bc_127) xor ad_127) xor ac_127);
    f_9(9) <= (((pkg_extract(f_8,9) xor bc_114) xor ad_114) xor ac_114);
    f_9(10) <= (((pkg_extract(f_8,10) xor bc_113) xor ad_113) xor ac_113);
    f_9(11) <= (((pkg_extract(f_8,11) xor bc_116) xor ad_116) xor ac_116);
    f_9(12) <= (((pkg_extract(f_8,12) xor bc_115) xor ad_115) xor ac_115);
  end process;

  process(e_9,bc_131,ad_131,bd_131,bc_130,ad_130,bd_130,bc_133,ad_133,bd_133,bc_132,ad_132,bd_132,bc_135,ad_135,bd_135,bc_134,ad_134,bd_134,bc_137,ad_137,bd_137,bc_136,ad_136,bd_136,bc_139,ad_139,bd_139,bc_138,ad_138,bd_138,bc_125,ad_125,bd_125,bc_129,ad_129,bd_129,bc_128,ad_128,bd_128)
  begin
    e_10(0) <= (((pkg_extract(e_9,0) xor bc_131) xor ad_131) xor bd_131);
    e_10(1) <= (((pkg_extract(e_9,1) xor bc_130) xor ad_130) xor bd_130);
    e_10(2) <= (((pkg_extract(e_9,2) xor bc_133) xor ad_133) xor bd_133);
    e_10(3) <= (((pkg_extract(e_9,3) xor bc_132) xor ad_132) xor bd_132);
    e_10(4) <= (((pkg_extract(e_9,4) xor bc_135) xor ad_135) xor bd_135);
    e_10(5) <= (((pkg_extract(e_9,5) xor bc_134) xor ad_134) xor bd_134);
    e_10(6) <= (((pkg_extract(e_9,6) xor bc_137) xor ad_137) xor bd_137);
    e_10(7) <= (((pkg_extract(e_9,7) xor bc_136) xor ad_136) xor bd_136);
    e_10(8) <= (((pkg_extract(e_9,8) xor bc_139) xor ad_139) xor bd_139);
    e_10(9) <= (((pkg_extract(e_9,9) xor bc_138) xor ad_138) xor bd_138);
    e_10(10) <= (((pkg_extract(e_9,10) xor bc_125) xor ad_125) xor bd_125);
    e_10(11) <= (((pkg_extract(e_9,11) xor bc_129) xor ad_129) xor bd_129);
    e_10(12) <= (((pkg_extract(e_9,12) xor bc_128) xor ad_128) xor bd_128);
  end process;

  process(f_9,bc_131,ad_131,ac_131,bc_130,ad_130,ac_130,bc_133,ad_133,ac_133,bc_132,ad_132,ac_132,bc_135,ad_135,ac_135,bc_134,ad_134,ac_134,bc_137,ad_137,ac_137,bc_136,ad_136,ac_136,bc_139,ad_139,ac_139,bc_138,ad_138,ac_138,bc_125,ad_125,ac_125,bc_129,ad_129,ac_129,bc_128,ad_128,ac_128)
  begin
    f_10(0) <= (((pkg_extract(f_9,0) xor bc_131) xor ad_131) xor ac_131);
    f_10(1) <= (((pkg_extract(f_9,1) xor bc_130) xor ad_130) xor ac_130);
    f_10(2) <= (((pkg_extract(f_9,2) xor bc_133) xor ad_133) xor ac_133);
    f_10(3) <= (((pkg_extract(f_9,3) xor bc_132) xor ad_132) xor ac_132);
    f_10(4) <= (((pkg_extract(f_9,4) xor bc_135) xor ad_135) xor ac_135);
    f_10(5) <= (((pkg_extract(f_9,5) xor bc_134) xor ad_134) xor ac_134);
    f_10(6) <= (((pkg_extract(f_9,6) xor bc_137) xor ad_137) xor ac_137);
    f_10(7) <= (((pkg_extract(f_9,7) xor bc_136) xor ad_136) xor ac_136);
    f_10(8) <= (((pkg_extract(f_9,8) xor bc_139) xor ad_139) xor ac_139);
    f_10(9) <= (((pkg_extract(f_9,9) xor bc_138) xor ad_138) xor ac_138);
    f_10(10) <= (((pkg_extract(f_9,10) xor bc_125) xor ad_125) xor ac_125);
    f_10(11) <= (((pkg_extract(f_9,11) xor bc_129) xor ad_129) xor ac_129);
    f_10(12) <= (((pkg_extract(f_9,12) xor bc_128) xor ad_128) xor ac_128);
  end process;

  process(e_10,bc_144,ad_144,bd_144,bc_143,ad_143,bd_143,bc_146,ad_146,bd_146,bc_145,ad_145,bd_145,bc_148,ad_148,bd_148,bc_147,ad_147,bd_147,bc_150,ad_150,bd_150,bc_149,ad_149,bd_149,bc_152,ad_152,bd_152,bc_151,ad_151,bd_151,bc_155,ad_155,bd_155,bc_142,ad_142,bd_142,bc_141,ad_141,bd_141)
  begin
    e_11(0) <= (((pkg_extract(e_10,0) xor bc_144) xor ad_144) xor bd_144);
    e_11(1) <= (((pkg_extract(e_10,1) xor bc_143) xor ad_143) xor bd_143);
    e_11(2) <= (((pkg_extract(e_10,2) xor bc_146) xor ad_146) xor bd_146);
    e_11(3) <= (((pkg_extract(e_10,3) xor bc_145) xor ad_145) xor bd_145);
    e_11(4) <= (((pkg_extract(e_10,4) xor bc_148) xor ad_148) xor bd_148);
    e_11(5) <= (((pkg_extract(e_10,5) xor bc_147) xor ad_147) xor bd_147);
    e_11(6) <= (((pkg_extract(e_10,6) xor bc_150) xor ad_150) xor bd_150);
    e_11(7) <= (((pkg_extract(e_10,7) xor bc_149) xor ad_149) xor bd_149);
    e_11(8) <= (((pkg_extract(e_10,8) xor bc_152) xor ad_152) xor bd_152);
    e_11(9) <= (((pkg_extract(e_10,9) xor bc_151) xor ad_151) xor bd_151);
    e_11(10) <= (((pkg_extract(e_10,10) xor bc_155) xor ad_155) xor bd_155);
    e_11(11) <= (((pkg_extract(e_10,11) xor bc_142) xor ad_142) xor bd_142);
    e_11(12) <= (((pkg_extract(e_10,12) xor bc_141) xor ad_141) xor bd_141);
  end process;

  process(f_10,bc_144,ad_144,ac_144,bc_143,ad_143,ac_143,bc_146,ad_146,ac_146,bc_145,ad_145,ac_145,bc_148,ad_148,ac_148,bc_147,ad_147,ac_147,bc_150,ad_150,ac_150,bc_149,ad_149,ac_149,bc_152,ad_152,ac_152,bc_151,ad_151,ac_151,bc_155,ad_155,ac_155,bc_142,ad_142,ac_142,bc_141,ad_141,ac_141)
  begin
    f_11(0) <= (((pkg_extract(f_10,0) xor bc_144) xor ad_144) xor ac_144);
    f_11(1) <= (((pkg_extract(f_10,1) xor bc_143) xor ad_143) xor ac_143);
    f_11(2) <= (((pkg_extract(f_10,2) xor bc_146) xor ad_146) xor ac_146);
    f_11(3) <= (((pkg_extract(f_10,3) xor bc_145) xor ad_145) xor ac_145);
    f_11(4) <= (((pkg_extract(f_10,4) xor bc_148) xor ad_148) xor ac_148);
    f_11(5) <= (((pkg_extract(f_10,5) xor bc_147) xor ad_147) xor ac_147);
    f_11(6) <= (((pkg_extract(f_10,6) xor bc_150) xor ad_150) xor ac_150);
    f_11(7) <= (((pkg_extract(f_10,7) xor bc_149) xor ad_149) xor ac_149);
    f_11(8) <= (((pkg_extract(f_10,8) xor bc_152) xor ad_152) xor ac_152);
    f_11(9) <= (((pkg_extract(f_10,9) xor bc_151) xor ad_151) xor ac_151);
    f_11(10) <= (((pkg_extract(f_10,10) xor bc_155) xor ad_155) xor ac_155);
    f_11(11) <= (((pkg_extract(f_10,11) xor bc_142) xor ad_142) xor ac_142);
    f_11(12) <= (((pkg_extract(f_10,12) xor bc_141) xor ad_141) xor ac_141);
  end process;

  process(e_11,bc_157,ad_157,bd_157,bc_156,ad_156,bd_156,bc_159,ad_159,bd_159,bc_158,ad_158,bd_158,bc_161,ad_161,bd_161,bc_160,ad_160,bd_160,bc_163,ad_163,bd_163,bc_162,ad_162,bd_162,bc_165,ad_165,bd_165,bc_164,ad_164,bd_164,bc_167,ad_167,bd_167,bc_166,ad_166,bd_166,bc_153,ad_153,bd_153)
  begin
    e_12(0) <= (((pkg_extract(e_11,0) xor bc_157) xor ad_157) xor bd_157);
    e_12(1) <= (((pkg_extract(e_11,1) xor bc_156) xor ad_156) xor bd_156);
    e_12(2) <= (((pkg_extract(e_11,2) xor bc_159) xor ad_159) xor bd_159);
    e_12(3) <= (((pkg_extract(e_11,3) xor bc_158) xor ad_158) xor bd_158);
    e_12(4) <= (((pkg_extract(e_11,4) xor bc_161) xor ad_161) xor bd_161);
    e_12(5) <= (((pkg_extract(e_11,5) xor bc_160) xor ad_160) xor bd_160);
    e_12(6) <= (((pkg_extract(e_11,6) xor bc_163) xor ad_163) xor bd_163);
    e_12(7) <= (((pkg_extract(e_11,7) xor bc_162) xor ad_162) xor bd_162);
    e_12(8) <= (((pkg_extract(e_11,8) xor bc_165) xor ad_165) xor bd_165);
    e_12(9) <= (((pkg_extract(e_11,9) xor bc_164) xor ad_164) xor bd_164);
    e_12(10) <= (((pkg_extract(e_11,10) xor bc_167) xor ad_167) xor bd_167);
    e_12(11) <= (((pkg_extract(e_11,11) xor bc_166) xor ad_166) xor bd_166);
    e_12(12) <= (((pkg_extract(e_11,12) xor bc_153) xor ad_153) xor bd_153);
  end process;

  process(f_11,bc_157,ad_157,ac_157,bc_156,ad_156,ac_156,bc_159,ad_159,ac_159,bc_158,ad_158,ac_158,bc_161,ad_161,ac_161,bc_160,ad_160,ac_160,bc_163,ad_163,ac_163,bc_162,ad_162,ac_162,bc_165,ad_165,ac_165,bc_164,ad_164,ac_164,bc_167,ad_167,ac_167,bc_166,ad_166,ac_166,bc_153,ad_153,ac_153)
  begin
    f_12(0) <= (((pkg_extract(f_11,0) xor bc_157) xor ad_157) xor ac_157);
    f_12(1) <= (((pkg_extract(f_11,1) xor bc_156) xor ad_156) xor ac_156);
    f_12(2) <= (((pkg_extract(f_11,2) xor bc_159) xor ad_159) xor ac_159);
    f_12(3) <= (((pkg_extract(f_11,3) xor bc_158) xor ad_158) xor ac_158);
    f_12(4) <= (((pkg_extract(f_11,4) xor bc_161) xor ad_161) xor ac_161);
    f_12(5) <= (((pkg_extract(f_11,5) xor bc_160) xor ad_160) xor ac_160);
    f_12(6) <= (((pkg_extract(f_11,6) xor bc_163) xor ad_163) xor ac_163);
    f_12(7) <= (((pkg_extract(f_11,7) xor bc_162) xor ad_162) xor ac_162);
    f_12(8) <= (((pkg_extract(f_11,8) xor bc_165) xor ad_165) xor ac_165);
    f_12(9) <= (((pkg_extract(f_11,9) xor bc_164) xor ad_164) xor ac_164);
    f_12(10) <= (((pkg_extract(f_11,10) xor bc_167) xor ad_167) xor ac_167);
    f_12(11) <= (((pkg_extract(f_11,11) xor bc_166) xor ad_166) xor ac_166);
    f_12(12) <= (((pkg_extract(f_11,12) xor bc_153) xor ad_153) xor ac_153);
  end process;

  io_z_0 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,0)),pkg_toStdLogicVector(pkg_extract(f_12,0)));
  io_z_1 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,1)),pkg_toStdLogicVector(pkg_extract(f_12,1)));
  io_z_2 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,2)),pkg_toStdLogicVector(pkg_extract(f_12,2)));
  io_z_3 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,3)),pkg_toStdLogicVector(pkg_extract(f_12,3)));
  io_z_4 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,4)),pkg_toStdLogicVector(pkg_extract(f_12,4)));
  io_z_5 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,5)),pkg_toStdLogicVector(pkg_extract(f_12,5)));
  io_z_6 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,6)),pkg_toStdLogicVector(pkg_extract(f_12,6)));
  io_z_7 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,7)),pkg_toStdLogicVector(pkg_extract(f_12,7)));
  io_z_8 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,8)),pkg_toStdLogicVector(pkg_extract(f_12,8)));
  io_z_9 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,9)),pkg_toStdLogicVector(pkg_extract(f_12,9)));
  io_z_10 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,10)),pkg_toStdLogicVector(pkg_extract(f_12,10)));
  io_z_11 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,11)),pkg_toStdLogicVector(pkg_extract(f_12,11)));
  io_z_12 <= pkg_cat(pkg_toStdLogicVector(pkg_extract(e_12,12)),pkg_toStdLogicVector(pkg_extract(f_12,12)));
end arch;


--G4MulTIMaskedN_1 replaced by G4MulTIMaskedN


--G4MulTIMaskedN_2 replaced by G4MulTIMaskedN

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity G4ScaleN is
  port(
    io_t : in std_logic_vector(1 downto 0);
    io_x : out std_logic_vector(1 downto 0)
  );
end G4ScaleN;

architecture arch of G4ScaleN is

begin
  io_x <= pkg_cat(pkg_toStdLogicVector(pkg_extract(io_t,0)),pkg_toStdLogicVector((pkg_extract(io_t,1) xor pkg_extract(io_t,0))));
end arch;


--G4ScaleN_1 replaced by G4ScaleN


--G4ScaleN_2 replaced by G4ScaleN


--G4ScaleN_3 replaced by G4ScaleN


--G4ScaleN_4 replaced by G4ScaleN


--G4ScaleN_5 replaced by G4ScaleN


--G4ScaleN_6 replaced by G4ScaleN


--G4ScaleN_7 replaced by G4ScaleN


--G4ScaleN_8 replaced by G4ScaleN


--G4ScaleN_9 replaced by G4ScaleN


--G4ScaleN_10 replaced by G4ScaleN


--G4ScaleN_11 replaced by G4ScaleN


--G4ScaleN_12 replaced by G4ScaleN


--G4MulTIMaskedN_3 replaced by G4MulTIMaskedN


--G4MulTIMaskedN_4 replaced by G4MulTIMaskedN


--G4MulTIMaskedN_5 replaced by G4MulTIMaskedN


--G4ScaleN_13 replaced by G4ScaleN


--G4ScaleN_14 replaced by G4ScaleN


--G4ScaleN_15 replaced by G4ScaleN


--G4ScaleN_16 replaced by G4ScaleN


--G4ScaleN_17 replaced by G4ScaleN


--G4ScaleN_18 replaced by G4ScaleN


--G4ScaleN_19 replaced by G4ScaleN


--G4ScaleN_20 replaced by G4ScaleN


--G4ScaleN_21 replaced by G4ScaleN


--G4ScaleN_22 replaced by G4ScaleN


--G4ScaleN_23 replaced by G4ScaleN


--G4ScaleN_24 replaced by G4ScaleN


--G4ScaleN_25 replaced by G4ScaleN


--G4MulTIMaskedN_6 replaced by G4MulTIMaskedN


--G4MulTIMaskedN_7 replaced by G4MulTIMaskedN


--G4MulTIMaskedN_8 replaced by G4MulTIMaskedN


--G4ScaleN_26 replaced by G4ScaleN


--G4ScaleN_27 replaced by G4ScaleN


--G4ScaleN_28 replaced by G4ScaleN


--G4ScaleN_29 replaced by G4ScaleN


--G4ScaleN_30 replaced by G4ScaleN


--G4ScaleN_31 replaced by G4ScaleN


--G4ScaleN_32 replaced by G4ScaleN


--G4ScaleN_33 replaced by G4ScaleN


--G4ScaleN_34 replaced by G4ScaleN


--G4ScaleN_35 replaced by G4ScaleN


--G4ScaleN_36 replaced by G4ScaleN


--G4ScaleN_37 replaced by G4ScaleN


--G4ScaleN_38 replaced by G4ScaleN


--G4MulTIMaskedN_9 replaced by G4MulTIMaskedN


--G4MulTIMaskedN_10 replaced by G4MulTIMaskedN


--G4MulTIMaskedN_11 replaced by G4MulTIMaskedN

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity G4Sq is
  port(
    io_t : in std_logic_vector(1 downto 0);
    io_x : out std_logic_vector(1 downto 0)
  );
end G4Sq;

architecture arch of G4Sq is

begin
  io_x <= pkg_cat(pkg_toStdLogicVector(pkg_extract(io_t,0)),pkg_toStdLogicVector(pkg_extract(io_t,1)));
end arch;


--G4ScaleN_39 replaced by G4ScaleN


--G4Sq_1 replaced by G4Sq


--G4ScaleN_40 replaced by G4ScaleN


--G4Sq_2 replaced by G4Sq


--G4ScaleN_41 replaced by G4ScaleN


--G4Sq_3 replaced by G4Sq


--G4ScaleN_42 replaced by G4ScaleN


--G4Sq_4 replaced by G4Sq


--G4ScaleN_43 replaced by G4ScaleN


--G4Sq_5 replaced by G4Sq


--G4ScaleN_44 replaced by G4ScaleN


--G4Sq_6 replaced by G4Sq


--G4ScaleN_45 replaced by G4ScaleN


--G4Sq_7 replaced by G4Sq


--G4ScaleN_46 replaced by G4ScaleN


--G4Sq_8 replaced by G4Sq


--G4ScaleN_47 replaced by G4ScaleN


--G4Sq_9 replaced by G4Sq


--G4ScaleN_48 replaced by G4ScaleN


--G4Sq_10 replaced by G4Sq


--G4ScaleN_49 replaced by G4ScaleN


--G4Sq_11 replaced by G4Sq


--G4ScaleN_50 replaced by G4ScaleN


--G4Sq_12 replaced by G4Sq


--G4ScaleN_51 replaced by G4ScaleN


--G4Sq_13 replaced by G4Sq


--G4Sq_14 replaced by G4Sq


--G4Sq_15 replaced by G4Sq


--G4Sq_16 replaced by G4Sq


--G4Sq_17 replaced by G4Sq


--G4Sq_18 replaced by G4Sq


--G4Sq_19 replaced by G4Sq


--G4Sq_20 replaced by G4Sq


--G4Sq_21 replaced by G4Sq


--G4Sq_22 replaced by G4Sq


--G4Sq_23 replaced by G4Sq


--G4Sq_24 replaced by G4Sq


--G4Sq_25 replaced by G4Sq


--G4Sq_26 replaced by G4Sq


--G4Sq_27 replaced by G4Sq

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity G4ScaleN2 is
  port(
    io_t : in std_logic_vector(1 downto 0);
    io_x : out std_logic_vector(1 downto 0)
  );
end G4ScaleN2;

architecture arch of G4ScaleN2 is

begin
  io_x <= pkg_cat(pkg_toStdLogicVector((pkg_extract(io_t,1) xor pkg_extract(io_t,0))),pkg_toStdLogicVector(pkg_extract(io_t,1)));
end arch;


--G4Sq_28 replaced by G4Sq


--G4Sq_29 replaced by G4Sq


--G4ScaleN2_1 replaced by G4ScaleN2


--G4Sq_30 replaced by G4Sq


--G4Sq_31 replaced by G4Sq


--G4ScaleN2_2 replaced by G4ScaleN2


--G4Sq_32 replaced by G4Sq


--G4Sq_33 replaced by G4Sq


--G4ScaleN2_3 replaced by G4ScaleN2


--G4Sq_34 replaced by G4Sq


--G4Sq_35 replaced by G4Sq


--G4ScaleN2_4 replaced by G4ScaleN2


--G4Sq_36 replaced by G4Sq


--G4Sq_37 replaced by G4Sq


--G4ScaleN2_5 replaced by G4ScaleN2


--G4Sq_38 replaced by G4Sq


--G4Sq_39 replaced by G4Sq


--G4ScaleN2_6 replaced by G4ScaleN2


--G4Sq_40 replaced by G4Sq


--G4Sq_41 replaced by G4Sq


--G4ScaleN2_7 replaced by G4ScaleN2


--G4Sq_42 replaced by G4Sq


--G4Sq_43 replaced by G4Sq


--G4ScaleN2_8 replaced by G4ScaleN2


--G4Sq_44 replaced by G4Sq


--G4Sq_45 replaced by G4Sq


--G4ScaleN2_9 replaced by G4ScaleN2


--G4Sq_46 replaced by G4Sq


--G4Sq_47 replaced by G4Sq


--G4ScaleN2_10 replaced by G4ScaleN2


--G4Sq_48 replaced by G4Sq


--G4Sq_49 replaced by G4Sq


--G4ScaleN2_11 replaced by G4ScaleN2


--G4Sq_50 replaced by G4Sq


--G4Sq_51 replaced by G4Sq


--G4ScaleN2_12 replaced by G4ScaleN2

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity G16MulTIMaskedN is
  port(
    io_x_0 : in std_logic_vector(3 downto 0);
    io_x_1 : in std_logic_vector(3 downto 0);
    io_x_2 : in std_logic_vector(3 downto 0);
    io_x_3 : in std_logic_vector(3 downto 0);
    io_x_4 : in std_logic_vector(3 downto 0);
    io_x_5 : in std_logic_vector(3 downto 0);
    io_x_6 : in std_logic_vector(3 downto 0);
    io_x_7 : in std_logic_vector(3 downto 0);
    io_x_8 : in std_logic_vector(3 downto 0);
    io_x_9 : in std_logic_vector(3 downto 0);
    io_x_10 : in std_logic_vector(3 downto 0);
    io_x_11 : in std_logic_vector(3 downto 0);
    io_x_12 : in std_logic_vector(3 downto 0);
    io_y_0 : in std_logic_vector(3 downto 0);
    io_y_1 : in std_logic_vector(3 downto 0);
    io_y_2 : in std_logic_vector(3 downto 0);
    io_y_3 : in std_logic_vector(3 downto 0);
    io_y_4 : in std_logic_vector(3 downto 0);
    io_y_5 : in std_logic_vector(3 downto 0);
    io_y_6 : in std_logic_vector(3 downto 0);
    io_y_7 : in std_logic_vector(3 downto 0);
    io_y_8 : in std_logic_vector(3 downto 0);
    io_y_9 : in std_logic_vector(3 downto 0);
    io_y_10 : in std_logic_vector(3 downto 0);
    io_y_11 : in std_logic_vector(3 downto 0);
    io_y_12 : in std_logic_vector(3 downto 0);
    io_z_0 : out std_logic_vector(3 downto 0);
    io_z_1 : out std_logic_vector(3 downto 0);
    io_z_2 : out std_logic_vector(3 downto 0);
    io_z_3 : out std_logic_vector(3 downto 0);
    io_z_4 : out std_logic_vector(3 downto 0);
    io_z_5 : out std_logic_vector(3 downto 0);
    io_z_6 : out std_logic_vector(3 downto 0);
    io_z_7 : out std_logic_vector(3 downto 0);
    io_z_8 : out std_logic_vector(3 downto 0);
    io_z_9 : out std_logic_vector(3 downto 0);
    io_z_10 : out std_logic_vector(3 downto 0);
    io_z_11 : out std_logic_vector(3 downto 0);
    io_z_12 : out std_logic_vector(3 downto 0);
    clk : in std_logic;
    reset : in std_logic
  );
end G16MulTIMaskedN;

architecture arch of G16MulTIMaskedN is
  signal mul1_io_x_0 : std_logic_vector(1 downto 0);
  signal mul1_io_x_1 : std_logic_vector(1 downto 0);
  signal mul1_io_x_2 : std_logic_vector(1 downto 0);
  signal mul1_io_x_3 : std_logic_vector(1 downto 0);
  signal mul1_io_x_4 : std_logic_vector(1 downto 0);
  signal mul1_io_x_5 : std_logic_vector(1 downto 0);
  signal mul1_io_x_6 : std_logic_vector(1 downto 0);
  signal mul1_io_x_7 : std_logic_vector(1 downto 0);
  signal mul1_io_x_8 : std_logic_vector(1 downto 0);
  signal mul1_io_x_9 : std_logic_vector(1 downto 0);
  signal mul1_io_x_10 : std_logic_vector(1 downto 0);
  signal mul1_io_x_11 : std_logic_vector(1 downto 0);
  signal mul1_io_x_12 : std_logic_vector(1 downto 0);
  signal mul1_io_y_0 : std_logic_vector(1 downto 0);
  signal mul1_io_y_1 : std_logic_vector(1 downto 0);
  signal mul1_io_y_2 : std_logic_vector(1 downto 0);
  signal mul1_io_y_3 : std_logic_vector(1 downto 0);
  signal mul1_io_y_4 : std_logic_vector(1 downto 0);
  signal mul1_io_y_5 : std_logic_vector(1 downto 0);
  signal mul1_io_y_6 : std_logic_vector(1 downto 0);
  signal mul1_io_y_7 : std_logic_vector(1 downto 0);
  signal mul1_io_y_8 : std_logic_vector(1 downto 0);
  signal mul1_io_y_9 : std_logic_vector(1 downto 0);
  signal mul1_io_y_10 : std_logic_vector(1 downto 0);
  signal mul1_io_y_11 : std_logic_vector(1 downto 0);
  signal mul1_io_y_12 : std_logic_vector(1 downto 0);
  signal mul1_io_z_0 : std_logic_vector(1 downto 0);
  signal mul1_io_z_1 : std_logic_vector(1 downto 0);
  signal mul1_io_z_2 : std_logic_vector(1 downto 0);
  signal mul1_io_z_3 : std_logic_vector(1 downto 0);
  signal mul1_io_z_4 : std_logic_vector(1 downto 0);
  signal mul1_io_z_5 : std_logic_vector(1 downto 0);
  signal mul1_io_z_6 : std_logic_vector(1 downto 0);
  signal mul1_io_z_7 : std_logic_vector(1 downto 0);
  signal mul1_io_z_8 : std_logic_vector(1 downto 0);
  signal mul1_io_z_9 : std_logic_vector(1 downto 0);
  signal mul1_io_z_10 : std_logic_vector(1 downto 0);
  signal mul1_io_z_11 : std_logic_vector(1 downto 0);
  signal mul1_io_z_12 : std_logic_vector(1 downto 0);
  signal mul2_io_z_0 : std_logic_vector(1 downto 0);
  signal mul2_io_z_1 : std_logic_vector(1 downto 0);
  signal mul2_io_z_2 : std_logic_vector(1 downto 0);
  signal mul2_io_z_3 : std_logic_vector(1 downto 0);
  signal mul2_io_z_4 : std_logic_vector(1 downto 0);
  signal mul2_io_z_5 : std_logic_vector(1 downto 0);
  signal mul2_io_z_6 : std_logic_vector(1 downto 0);
  signal mul2_io_z_7 : std_logic_vector(1 downto 0);
  signal mul2_io_z_8 : std_logic_vector(1 downto 0);
  signal mul2_io_z_9 : std_logic_vector(1 downto 0);
  signal mul2_io_z_10 : std_logic_vector(1 downto 0);
  signal mul2_io_z_11 : std_logic_vector(1 downto 0);
  signal mul2_io_z_12 : std_logic_vector(1 downto 0);
  signal mul3_io_z_0 : std_logic_vector(1 downto 0);
  signal mul3_io_z_1 : std_logic_vector(1 downto 0);
  signal mul3_io_z_2 : std_logic_vector(1 downto 0);
  signal mul3_io_z_3 : std_logic_vector(1 downto 0);
  signal mul3_io_z_4 : std_logic_vector(1 downto 0);
  signal mul3_io_z_5 : std_logic_vector(1 downto 0);
  signal mul3_io_z_6 : std_logic_vector(1 downto 0);
  signal mul3_io_z_7 : std_logic_vector(1 downto 0);
  signal mul3_io_z_8 : std_logic_vector(1 downto 0);
  signal mul3_io_z_9 : std_logic_vector(1 downto 0);
  signal mul3_io_z_10 : std_logic_vector(1 downto 0);
  signal mul3_io_z_11 : std_logic_vector(1 downto 0);
  signal mul3_io_z_12 : std_logic_vector(1 downto 0);
  signal g4ScaleN_52_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_53_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_54_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_55_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_56_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_57_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_58_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_59_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_60_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_61_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_62_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_63_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_64_io_x : std_logic_vector(1 downto 0);

  signal dummy : std_logic;
  signal a_0 : std_logic_vector(1 downto 0);
  signal a_1 : std_logic_vector(1 downto 0);
  signal a_2 : std_logic_vector(1 downto 0);
  signal a_3 : std_logic_vector(1 downto 0);
  signal a_4 : std_logic_vector(1 downto 0);
  signal a_5 : std_logic_vector(1 downto 0);
  signal a_6 : std_logic_vector(1 downto 0);
  signal a_7 : std_logic_vector(1 downto 0);
  signal a_8 : std_logic_vector(1 downto 0);
  signal a_9 : std_logic_vector(1 downto 0);
  signal a_10 : std_logic_vector(1 downto 0);
  signal a_11 : std_logic_vector(1 downto 0);
  signal a_12 : std_logic_vector(1 downto 0);
  signal b_0 : std_logic_vector(1 downto 0);
  signal b_1 : std_logic_vector(1 downto 0);
  signal b_2 : std_logic_vector(1 downto 0);
  signal b_3 : std_logic_vector(1 downto 0);
  signal b_4 : std_logic_vector(1 downto 0);
  signal b_5 : std_logic_vector(1 downto 0);
  signal b_6 : std_logic_vector(1 downto 0);
  signal b_7 : std_logic_vector(1 downto 0);
  signal b_8 : std_logic_vector(1 downto 0);
  signal b_9 : std_logic_vector(1 downto 0);
  signal b_10 : std_logic_vector(1 downto 0);
  signal b_11 : std_logic_vector(1 downto 0);
  signal b_12 : std_logic_vector(1 downto 0);
  signal c_0 : std_logic_vector(1 downto 0);
  signal c_1 : std_logic_vector(1 downto 0);
  signal c_2 : std_logic_vector(1 downto 0);
  signal c_3 : std_logic_vector(1 downto 0);
  signal c_4 : std_logic_vector(1 downto 0);
  signal c_5 : std_logic_vector(1 downto 0);
  signal c_6 : std_logic_vector(1 downto 0);
  signal c_7 : std_logic_vector(1 downto 0);
  signal c_8 : std_logic_vector(1 downto 0);
  signal c_9 : std_logic_vector(1 downto 0);
  signal c_10 : std_logic_vector(1 downto 0);
  signal c_11 : std_logic_vector(1 downto 0);
  signal c_12 : std_logic_vector(1 downto 0);
  signal d_0 : std_logic_vector(1 downto 0);
  signal d_1 : std_logic_vector(1 downto 0);
  signal d_2 : std_logic_vector(1 downto 0);
  signal d_3 : std_logic_vector(1 downto 0);
  signal d_4 : std_logic_vector(1 downto 0);
  signal d_5 : std_logic_vector(1 downto 0);
  signal d_6 : std_logic_vector(1 downto 0);
  signal d_7 : std_logic_vector(1 downto 0);
  signal d_8 : std_logic_vector(1 downto 0);
  signal d_9 : std_logic_vector(1 downto 0);
  signal d_10 : std_logic_vector(1 downto 0);
  signal d_11 : std_logic_vector(1 downto 0);
  signal d_12 : std_logic_vector(1 downto 0);
  signal e_0 : std_logic_vector(1 downto 0);
  signal e_1 : std_logic_vector(1 downto 0);
  signal e_2 : std_logic_vector(1 downto 0);
  signal e_3 : std_logic_vector(1 downto 0);
  signal e_4 : std_logic_vector(1 downto 0);
  signal e_5 : std_logic_vector(1 downto 0);
  signal e_6 : std_logic_vector(1 downto 0);
  signal e_7 : std_logic_vector(1 downto 0);
  signal e_8 : std_logic_vector(1 downto 0);
  signal e_9 : std_logic_vector(1 downto 0);
  signal e_10 : std_logic_vector(1 downto 0);
  signal e_11 : std_logic_vector(1 downto 0);
  signal e_12 : std_logic_vector(1 downto 0);
  signal f_0 : std_logic_vector(1 downto 0);
  signal f_1 : std_logic_vector(1 downto 0);
  signal f_2 : std_logic_vector(1 downto 0);
  signal f_3 : std_logic_vector(1 downto 0);
  signal f_4 : std_logic_vector(1 downto 0);
  signal f_5 : std_logic_vector(1 downto 0);
  signal f_6 : std_logic_vector(1 downto 0);
  signal f_7 : std_logic_vector(1 downto 0);
  signal f_8 : std_logic_vector(1 downto 0);
  signal f_9 : std_logic_vector(1 downto 0);
  signal f_10 : std_logic_vector(1 downto 0);
  signal f_11 : std_logic_vector(1 downto 0);
  signal f_12 : std_logic_vector(1 downto 0);
  signal g_0 : std_logic_vector(1 downto 0);
  signal g_1 : std_logic_vector(1 downto 0);
  signal g_2 : std_logic_vector(1 downto 0);
  signal g_3 : std_logic_vector(1 downto 0);
  signal g_4 : std_logic_vector(1 downto 0);
  signal g_5 : std_logic_vector(1 downto 0);
  signal g_6 : std_logic_vector(1 downto 0);
  signal g_7 : std_logic_vector(1 downto 0);
  signal g_8 : std_logic_vector(1 downto 0);
  signal g_9 : std_logic_vector(1 downto 0);
  signal g_10 : std_logic_vector(1 downto 0);
  signal g_11 : std_logic_vector(1 downto 0);
  signal g_12 : std_logic_vector(1 downto 0);
  signal h_0 : std_logic_vector(1 downto 0);
  signal h_1 : std_logic_vector(1 downto 0);
  signal h_2 : std_logic_vector(1 downto 0);
  signal h_3 : std_logic_vector(1 downto 0);
  signal h_4 : std_logic_vector(1 downto 0);
  signal h_5 : std_logic_vector(1 downto 0);
  signal h_6 : std_logic_vector(1 downto 0);
  signal h_7 : std_logic_vector(1 downto 0);
  signal h_8 : std_logic_vector(1 downto 0);
  signal h_9 : std_logic_vector(1 downto 0);
  signal h_10 : std_logic_vector(1 downto 0);
  signal h_11 : std_logic_vector(1 downto 0);
  signal h_12 : std_logic_vector(1 downto 0);
  signal p_0 : std_logic_vector(1 downto 0);
  signal p_1 : std_logic_vector(1 downto 0);
  signal p_2 : std_logic_vector(1 downto 0);
  signal p_3 : std_logic_vector(1 downto 0);
  signal p_4 : std_logic_vector(1 downto 0);
  signal p_5 : std_logic_vector(1 downto 0);
  signal p_6 : std_logic_vector(1 downto 0);
  signal p_7 : std_logic_vector(1 downto 0);
  signal p_8 : std_logic_vector(1 downto 0);
  signal p_9 : std_logic_vector(1 downto 0);
  signal p_10 : std_logic_vector(1 downto 0);
  signal p_11 : std_logic_vector(1 downto 0);
  signal p_12 : std_logic_vector(1 downto 0);
  signal q_0 : std_logic_vector(1 downto 0);
  signal q_1 : std_logic_vector(1 downto 0);
  signal q_2 : std_logic_vector(1 downto 0);
  signal q_3 : std_logic_vector(1 downto 0);
  signal q_4 : std_logic_vector(1 downto 0);
  signal q_5 : std_logic_vector(1 downto 0);
  signal q_6 : std_logic_vector(1 downto 0);
  signal q_7 : std_logic_vector(1 downto 0);
  signal q_8 : std_logic_vector(1 downto 0);
  signal q_9 : std_logic_vector(1 downto 0);
  signal q_10 : std_logic_vector(1 downto 0);
  signal q_11 : std_logic_vector(1 downto 0);
  signal q_12 : std_logic_vector(1 downto 0);
begin
  mul1 : entity work.G4MulTIMaskedN
    port map ( 
      io_x_0 => mul1_io_x_0,
      io_x_1 => mul1_io_x_1,
      io_x_2 => mul1_io_x_2,
      io_x_3 => mul1_io_x_3,
      io_x_4 => mul1_io_x_4,
      io_x_5 => mul1_io_x_5,
      io_x_6 => mul1_io_x_6,
      io_x_7 => mul1_io_x_7,
      io_x_8 => mul1_io_x_8,
      io_x_9 => mul1_io_x_9,
      io_x_10 => mul1_io_x_10,
      io_x_11 => mul1_io_x_11,
      io_x_12 => mul1_io_x_12,
      io_y_0 => mul1_io_y_0,
      io_y_1 => mul1_io_y_1,
      io_y_2 => mul1_io_y_2,
      io_y_3 => mul1_io_y_3,
      io_y_4 => mul1_io_y_4,
      io_y_5 => mul1_io_y_5,
      io_y_6 => mul1_io_y_6,
      io_y_7 => mul1_io_y_7,
      io_y_8 => mul1_io_y_8,
      io_y_9 => mul1_io_y_9,
      io_y_10 => mul1_io_y_10,
      io_y_11 => mul1_io_y_11,
      io_y_12 => mul1_io_y_12,
      io_z_0 => mul1_io_z_0,
      io_z_1 => mul1_io_z_1,
      io_z_2 => mul1_io_z_2,
      io_z_3 => mul1_io_z_3,
      io_z_4 => mul1_io_z_4,
      io_z_5 => mul1_io_z_5,
      io_z_6 => mul1_io_z_6,
      io_z_7 => mul1_io_z_7,
      io_z_8 => mul1_io_z_8,
      io_z_9 => mul1_io_z_9,
      io_z_10 => mul1_io_z_10,
      io_z_11 => mul1_io_z_11,
      io_z_12 => mul1_io_z_12,
      clk => clk,
      reset => reset 
    );
  mul2 : entity work.G4MulTIMaskedN
    port map ( 
      io_x_0 => a_0,
      io_x_1 => a_1,
      io_x_2 => a_2,
      io_x_3 => a_3,
      io_x_4 => a_4,
      io_x_5 => a_5,
      io_x_6 => a_6,
      io_x_7 => a_7,
      io_x_8 => a_8,
      io_x_9 => a_9,
      io_x_10 => a_10,
      io_x_11 => a_11,
      io_x_12 => a_12,
      io_y_0 => c_0,
      io_y_1 => c_1,
      io_y_2 => c_2,
      io_y_3 => c_3,
      io_y_4 => c_4,
      io_y_5 => c_5,
      io_y_6 => c_6,
      io_y_7 => c_7,
      io_y_8 => c_8,
      io_y_9 => c_9,
      io_y_10 => c_10,
      io_y_11 => c_11,
      io_y_12 => c_12,
      io_z_0 => mul2_io_z_0,
      io_z_1 => mul2_io_z_1,
      io_z_2 => mul2_io_z_2,
      io_z_3 => mul2_io_z_3,
      io_z_4 => mul2_io_z_4,
      io_z_5 => mul2_io_z_5,
      io_z_6 => mul2_io_z_6,
      io_z_7 => mul2_io_z_7,
      io_z_8 => mul2_io_z_8,
      io_z_9 => mul2_io_z_9,
      io_z_10 => mul2_io_z_10,
      io_z_11 => mul2_io_z_11,
      io_z_12 => mul2_io_z_12,
      clk => clk,
      reset => reset 
    );
  mul3 : entity work.G4MulTIMaskedN
    port map ( 
      io_x_0 => b_0,
      io_x_1 => b_1,
      io_x_2 => b_2,
      io_x_3 => b_3,
      io_x_4 => b_4,
      io_x_5 => b_5,
      io_x_6 => b_6,
      io_x_7 => b_7,
      io_x_8 => b_8,
      io_x_9 => b_9,
      io_x_10 => b_10,
      io_x_11 => b_11,
      io_x_12 => b_12,
      io_y_0 => d_0,
      io_y_1 => d_1,
      io_y_2 => d_2,
      io_y_3 => d_3,
      io_y_4 => d_4,
      io_y_5 => d_5,
      io_y_6 => d_6,
      io_y_7 => d_7,
      io_y_8 => d_8,
      io_y_9 => d_9,
      io_y_10 => d_10,
      io_y_11 => d_11,
      io_y_12 => d_12,
      io_z_0 => mul3_io_z_0,
      io_z_1 => mul3_io_z_1,
      io_z_2 => mul3_io_z_2,
      io_z_3 => mul3_io_z_3,
      io_z_4 => mul3_io_z_4,
      io_z_5 => mul3_io_z_5,
      io_z_6 => mul3_io_z_6,
      io_z_7 => mul3_io_z_7,
      io_z_8 => mul3_io_z_8,
      io_z_9 => mul3_io_z_9,
      io_z_10 => mul3_io_z_10,
      io_z_11 => mul3_io_z_11,
      io_z_12 => mul3_io_z_12,
      clk => clk,
      reset => reset 
    );
  g4ScaleN_52 : entity work.G4ScaleN
    port map ( 
      io_t => e_0,
      io_x => g4ScaleN_52_io_x 
    );
  g4ScaleN_53 : entity work.G4ScaleN
    port map ( 
      io_t => e_1,
      io_x => g4ScaleN_53_io_x 
    );
  g4ScaleN_54 : entity work.G4ScaleN
    port map ( 
      io_t => e_2,
      io_x => g4ScaleN_54_io_x 
    );
  g4ScaleN_55 : entity work.G4ScaleN
    port map ( 
      io_t => e_3,
      io_x => g4ScaleN_55_io_x 
    );
  g4ScaleN_56 : entity work.G4ScaleN
    port map ( 
      io_t => e_4,
      io_x => g4ScaleN_56_io_x 
    );
  g4ScaleN_57 : entity work.G4ScaleN
    port map ( 
      io_t => e_5,
      io_x => g4ScaleN_57_io_x 
    );
  g4ScaleN_58 : entity work.G4ScaleN
    port map ( 
      io_t => e_6,
      io_x => g4ScaleN_58_io_x 
    );
  g4ScaleN_59 : entity work.G4ScaleN
    port map ( 
      io_t => e_7,
      io_x => g4ScaleN_59_io_x 
    );
  g4ScaleN_60 : entity work.G4ScaleN
    port map ( 
      io_t => e_8,
      io_x => g4ScaleN_60_io_x 
    );
  g4ScaleN_61 : entity work.G4ScaleN
    port map ( 
      io_t => e_9,
      io_x => g4ScaleN_61_io_x 
    );
  g4ScaleN_62 : entity work.G4ScaleN
    port map ( 
      io_t => e_10,
      io_x => g4ScaleN_62_io_x 
    );
  g4ScaleN_63 : entity work.G4ScaleN
    port map ( 
      io_t => e_11,
      io_x => g4ScaleN_63_io_x 
    );
  g4ScaleN_64 : entity work.G4ScaleN
    port map ( 
      io_t => e_12,
      io_x => g4ScaleN_64_io_x 
    );
  dummy <= pkg_toStdLogic(false);
  a_0 <= pkg_extract(io_x_0,3,2);
  b_0 <= pkg_extract(io_x_0,1,0);
  c_0 <= pkg_extract(io_y_0,3,2);
  d_0 <= pkg_extract(io_y_0,1,0);
  a_1 <= pkg_extract(io_x_1,3,2);
  b_1 <= pkg_extract(io_x_1,1,0);
  c_1 <= pkg_extract(io_y_1,3,2);
  d_1 <= pkg_extract(io_y_1,1,0);
  a_2 <= pkg_extract(io_x_2,3,2);
  b_2 <= pkg_extract(io_x_2,1,0);
  c_2 <= pkg_extract(io_y_2,3,2);
  d_2 <= pkg_extract(io_y_2,1,0);
  a_3 <= pkg_extract(io_x_3,3,2);
  b_3 <= pkg_extract(io_x_3,1,0);
  c_3 <= pkg_extract(io_y_3,3,2);
  d_3 <= pkg_extract(io_y_3,1,0);
  a_4 <= pkg_extract(io_x_4,3,2);
  b_4 <= pkg_extract(io_x_4,1,0);
  c_4 <= pkg_extract(io_y_4,3,2);
  d_4 <= pkg_extract(io_y_4,1,0);
  a_5 <= pkg_extract(io_x_5,3,2);
  b_5 <= pkg_extract(io_x_5,1,0);
  c_5 <= pkg_extract(io_y_5,3,2);
  d_5 <= pkg_extract(io_y_5,1,0);
  a_6 <= pkg_extract(io_x_6,3,2);
  b_6 <= pkg_extract(io_x_6,1,0);
  c_6 <= pkg_extract(io_y_6,3,2);
  d_6 <= pkg_extract(io_y_6,1,0);
  a_7 <= pkg_extract(io_x_7,3,2);
  b_7 <= pkg_extract(io_x_7,1,0);
  c_7 <= pkg_extract(io_y_7,3,2);
  d_7 <= pkg_extract(io_y_7,1,0);
  a_8 <= pkg_extract(io_x_8,3,2);
  b_8 <= pkg_extract(io_x_8,1,0);
  c_8 <= pkg_extract(io_y_8,3,2);
  d_8 <= pkg_extract(io_y_8,1,0);
  a_9 <= pkg_extract(io_x_9,3,2);
  b_9 <= pkg_extract(io_x_9,1,0);
  c_9 <= pkg_extract(io_y_9,3,2);
  d_9 <= pkg_extract(io_y_9,1,0);
  a_10 <= pkg_extract(io_x_10,3,2);
  b_10 <= pkg_extract(io_x_10,1,0);
  c_10 <= pkg_extract(io_y_10,3,2);
  d_10 <= pkg_extract(io_y_10,1,0);
  a_11 <= pkg_extract(io_x_11,3,2);
  b_11 <= pkg_extract(io_x_11,1,0);
  c_11 <= pkg_extract(io_y_11,3,2);
  d_11 <= pkg_extract(io_y_11,1,0);
  a_12 <= pkg_extract(io_x_12,3,2);
  b_12 <= pkg_extract(io_x_12,1,0);
  c_12 <= pkg_extract(io_y_12,3,2);
  d_12 <= pkg_extract(io_y_12,1,0);
  mul1_io_x_0 <= (a_0 xor b_0);
  mul1_io_x_1 <= (a_1 xor b_1);
  mul1_io_x_2 <= (a_2 xor b_2);
  mul1_io_x_3 <= (a_3 xor b_3);
  mul1_io_x_4 <= (a_4 xor b_4);
  mul1_io_x_5 <= (a_5 xor b_5);
  mul1_io_x_6 <= (a_6 xor b_6);
  mul1_io_x_7 <= (a_7 xor b_7);
  mul1_io_x_8 <= (a_8 xor b_8);
  mul1_io_x_9 <= (a_9 xor b_9);
  mul1_io_x_10 <= (a_10 xor b_10);
  mul1_io_x_11 <= (a_11 xor b_11);
  mul1_io_x_12 <= (a_12 xor b_12);
  mul1_io_y_0 <= (c_0 xor d_0);
  mul1_io_y_1 <= (c_1 xor d_1);
  mul1_io_y_2 <= (c_2 xor d_2);
  mul1_io_y_3 <= (c_3 xor d_3);
  mul1_io_y_4 <= (c_4 xor d_4);
  mul1_io_y_5 <= (c_5 xor d_5);
  mul1_io_y_6 <= (c_6 xor d_6);
  mul1_io_y_7 <= (c_7 xor d_7);
  mul1_io_y_8 <= (c_8 xor d_8);
  mul1_io_y_9 <= (c_9 xor d_9);
  mul1_io_y_10 <= (c_10 xor d_10);
  mul1_io_y_11 <= (c_11 xor d_11);
  mul1_io_y_12 <= (c_12 xor d_12);
  e_0 <= mul1_io_z_0;
  e_1 <= mul1_io_z_1;
  e_2 <= mul1_io_z_2;
  e_3 <= mul1_io_z_3;
  e_4 <= mul1_io_z_4;
  e_5 <= mul1_io_z_5;
  e_6 <= mul1_io_z_6;
  e_7 <= mul1_io_z_7;
  e_8 <= mul1_io_z_8;
  e_9 <= mul1_io_z_9;
  e_10 <= mul1_io_z_10;
  e_11 <= mul1_io_z_11;
  e_12 <= mul1_io_z_12;
  f_0 <= g4ScaleN_52_io_x;
  f_1 <= g4ScaleN_53_io_x;
  f_2 <= g4ScaleN_54_io_x;
  f_3 <= g4ScaleN_55_io_x;
  f_4 <= g4ScaleN_56_io_x;
  f_5 <= g4ScaleN_57_io_x;
  f_6 <= g4ScaleN_58_io_x;
  f_7 <= g4ScaleN_59_io_x;
  f_8 <= g4ScaleN_60_io_x;
  f_9 <= g4ScaleN_61_io_x;
  f_10 <= g4ScaleN_62_io_x;
  f_11 <= g4ScaleN_63_io_x;
  f_12 <= g4ScaleN_64_io_x;
  g_0 <= mul2_io_z_0;
  g_1 <= mul2_io_z_1;
  g_2 <= mul2_io_z_2;
  g_3 <= mul2_io_z_3;
  g_4 <= mul2_io_z_4;
  g_5 <= mul2_io_z_5;
  g_6 <= mul2_io_z_6;
  g_7 <= mul2_io_z_7;
  g_8 <= mul2_io_z_8;
  g_9 <= mul2_io_z_9;
  g_10 <= mul2_io_z_10;
  g_11 <= mul2_io_z_11;
  g_12 <= mul2_io_z_12;
  h_0 <= mul3_io_z_0;
  h_1 <= mul3_io_z_1;
  h_2 <= mul3_io_z_2;
  h_3 <= mul3_io_z_3;
  h_4 <= mul3_io_z_4;
  h_5 <= mul3_io_z_5;
  h_6 <= mul3_io_z_6;
  h_7 <= mul3_io_z_7;
  h_8 <= mul3_io_z_8;
  h_9 <= mul3_io_z_9;
  h_10 <= mul3_io_z_10;
  h_11 <= mul3_io_z_11;
  h_12 <= mul3_io_z_12;
  p_0 <= (f_0 xor g_0);
  p_1 <= (f_1 xor g_1);
  p_2 <= (f_2 xor g_2);
  p_3 <= (f_3 xor g_3);
  p_4 <= (f_4 xor g_4);
  p_5 <= (f_5 xor g_5);
  p_6 <= (f_6 xor g_6);
  p_7 <= (f_7 xor g_7);
  p_8 <= (f_8 xor g_8);
  p_9 <= (f_9 xor g_9);
  p_10 <= (f_10 xor g_10);
  p_11 <= (f_11 xor g_11);
  p_12 <= (f_12 xor g_12);
  q_0 <= (f_0 xor h_0);
  q_1 <= (f_1 xor h_1);
  q_2 <= (f_2 xor h_2);
  q_3 <= (f_3 xor h_3);
  q_4 <= (f_4 xor h_4);
  q_5 <= (f_5 xor h_5);
  q_6 <= (f_6 xor h_6);
  q_7 <= (f_7 xor h_7);
  q_8 <= (f_8 xor h_8);
  q_9 <= (f_9 xor h_9);
  q_10 <= (f_10 xor h_10);
  q_11 <= (f_11 xor h_11);
  q_12 <= (f_12 xor h_12);
  io_z_0 <= pkg_cat(p_0,q_0);
  io_z_1 <= pkg_cat(p_1,q_1);
  io_z_2 <= pkg_cat(p_2,q_2);
  io_z_3 <= pkg_cat(p_3,q_3);
  io_z_4 <= pkg_cat(p_4,q_4);
  io_z_5 <= pkg_cat(p_5,q_5);
  io_z_6 <= pkg_cat(p_6,q_6);
  io_z_7 <= pkg_cat(p_7,q_7);
  io_z_8 <= pkg_cat(p_8,q_8);
  io_z_9 <= pkg_cat(p_9,q_9);
  io_z_10 <= pkg_cat(p_10,q_10);
  io_z_11 <= pkg_cat(p_11,q_11);
  io_z_12 <= pkg_cat(p_12,q_12);
end arch;


--G16MulTIMaskedN_1 replaced by G16MulTIMaskedN


--G16MulTIMaskedN_2 replaced by G16MulTIMaskedN

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity G16InvTIMaskedN is
  port(
    io_x_0 : in std_logic_vector(3 downto 0);
    io_x_1 : in std_logic_vector(3 downto 0);
    io_x_2 : in std_logic_vector(3 downto 0);
    io_x_3 : in std_logic_vector(3 downto 0);
    io_x_4 : in std_logic_vector(3 downto 0);
    io_x_5 : in std_logic_vector(3 downto 0);
    io_x_6 : in std_logic_vector(3 downto 0);
    io_x_7 : in std_logic_vector(3 downto 0);
    io_x_8 : in std_logic_vector(3 downto 0);
    io_x_9 : in std_logic_vector(3 downto 0);
    io_x_10 : in std_logic_vector(3 downto 0);
    io_x_11 : in std_logic_vector(3 downto 0);
    io_x_12 : in std_logic_vector(3 downto 0);
    io_z_0 : out std_logic_vector(3 downto 0);
    io_z_1 : out std_logic_vector(3 downto 0);
    io_z_2 : out std_logic_vector(3 downto 0);
    io_z_3 : out std_logic_vector(3 downto 0);
    io_z_4 : out std_logic_vector(3 downto 0);
    io_z_5 : out std_logic_vector(3 downto 0);
    io_z_6 : out std_logic_vector(3 downto 0);
    io_z_7 : out std_logic_vector(3 downto 0);
    io_z_8 : out std_logic_vector(3 downto 0);
    io_z_9 : out std_logic_vector(3 downto 0);
    io_z_10 : out std_logic_vector(3 downto 0);
    io_z_11 : out std_logic_vector(3 downto 0);
    io_z_12 : out std_logic_vector(3 downto 0);
    clk : in std_logic;
    reset : in std_logic
  );
end G16InvTIMaskedN;

architecture arch of G16InvTIMaskedN is
  signal g4Sq_65_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_66_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_67_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_68_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_69_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_70_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_71_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_72_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_73_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_74_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_75_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_76_io_t : std_logic_vector(1 downto 0);
  signal g4Sq_77_io_t : std_logic_vector(1 downto 0);
  signal mul1_io_z_0 : std_logic_vector(1 downto 0);
  signal mul1_io_z_1 : std_logic_vector(1 downto 0);
  signal mul1_io_z_2 : std_logic_vector(1 downto 0);
  signal mul1_io_z_3 : std_logic_vector(1 downto 0);
  signal mul1_io_z_4 : std_logic_vector(1 downto 0);
  signal mul1_io_z_5 : std_logic_vector(1 downto 0);
  signal mul1_io_z_6 : std_logic_vector(1 downto 0);
  signal mul1_io_z_7 : std_logic_vector(1 downto 0);
  signal mul1_io_z_8 : std_logic_vector(1 downto 0);
  signal mul1_io_z_9 : std_logic_vector(1 downto 0);
  signal mul1_io_z_10 : std_logic_vector(1 downto 0);
  signal mul1_io_z_11 : std_logic_vector(1 downto 0);
  signal mul1_io_z_12 : std_logic_vector(1 downto 0);
  signal mul2_io_z_0 : std_logic_vector(1 downto 0);
  signal mul2_io_z_1 : std_logic_vector(1 downto 0);
  signal mul2_io_z_2 : std_logic_vector(1 downto 0);
  signal mul2_io_z_3 : std_logic_vector(1 downto 0);
  signal mul2_io_z_4 : std_logic_vector(1 downto 0);
  signal mul2_io_z_5 : std_logic_vector(1 downto 0);
  signal mul2_io_z_6 : std_logic_vector(1 downto 0);
  signal mul2_io_z_7 : std_logic_vector(1 downto 0);
  signal mul2_io_z_8 : std_logic_vector(1 downto 0);
  signal mul2_io_z_9 : std_logic_vector(1 downto 0);
  signal mul2_io_z_10 : std_logic_vector(1 downto 0);
  signal mul2_io_z_11 : std_logic_vector(1 downto 0);
  signal mul2_io_z_12 : std_logic_vector(1 downto 0);
  signal mul3_io_z_0 : std_logic_vector(1 downto 0);
  signal mul3_io_z_1 : std_logic_vector(1 downto 0);
  signal mul3_io_z_2 : std_logic_vector(1 downto 0);
  signal mul3_io_z_3 : std_logic_vector(1 downto 0);
  signal mul3_io_z_4 : std_logic_vector(1 downto 0);
  signal mul3_io_z_5 : std_logic_vector(1 downto 0);
  signal mul3_io_z_6 : std_logic_vector(1 downto 0);
  signal mul3_io_z_7 : std_logic_vector(1 downto 0);
  signal mul3_io_z_8 : std_logic_vector(1 downto 0);
  signal mul3_io_z_9 : std_logic_vector(1 downto 0);
  signal mul3_io_z_10 : std_logic_vector(1 downto 0);
  signal mul3_io_z_11 : std_logic_vector(1 downto 0);
  signal mul3_io_z_12 : std_logic_vector(1 downto 0);
  signal g4Sq_52_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_52_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_53_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_53_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_54_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_54_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_55_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_55_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_56_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_56_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_57_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_57_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_58_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_58_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_59_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_59_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_60_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_60_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_61_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_61_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_62_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_62_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_63_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_63_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_64_io_x : std_logic_vector(1 downto 0);
  signal g4ScaleN_64_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_65_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_66_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_67_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_68_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_69_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_70_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_71_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_72_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_73_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_74_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_75_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_76_io_x : std_logic_vector(1 downto 0);
  signal g4Sq_77_io_x : std_logic_vector(1 downto 0);

  signal dummy : std_logic;
  signal a_0 : std_logic_vector(1 downto 0);
  signal a_1 : std_logic_vector(1 downto 0);
  signal a_2 : std_logic_vector(1 downto 0);
  signal a_3 : std_logic_vector(1 downto 0);
  signal a_4 : std_logic_vector(1 downto 0);
  signal a_5 : std_logic_vector(1 downto 0);
  signal a_6 : std_logic_vector(1 downto 0);
  signal a_7 : std_logic_vector(1 downto 0);
  signal a_8 : std_logic_vector(1 downto 0);
  signal a_9 : std_logic_vector(1 downto 0);
  signal a_10 : std_logic_vector(1 downto 0);
  signal a_11 : std_logic_vector(1 downto 0);
  signal a_12 : std_logic_vector(1 downto 0);
  signal b_0 : std_logic_vector(1 downto 0);
  signal b_1 : std_logic_vector(1 downto 0);
  signal b_2 : std_logic_vector(1 downto 0);
  signal b_3 : std_logic_vector(1 downto 0);
  signal b_4 : std_logic_vector(1 downto 0);
  signal b_5 : std_logic_vector(1 downto 0);
  signal b_6 : std_logic_vector(1 downto 0);
  signal b_7 : std_logic_vector(1 downto 0);
  signal b_8 : std_logic_vector(1 downto 0);
  signal b_9 : std_logic_vector(1 downto 0);
  signal b_10 : std_logic_vector(1 downto 0);
  signal b_11 : std_logic_vector(1 downto 0);
  signal b_12 : std_logic_vector(1 downto 0);
  signal c_0 : std_logic_vector(1 downto 0);
  signal c_1 : std_logic_vector(1 downto 0);
  signal c_2 : std_logic_vector(1 downto 0);
  signal c_3 : std_logic_vector(1 downto 0);
  signal c_4 : std_logic_vector(1 downto 0);
  signal c_5 : std_logic_vector(1 downto 0);
  signal c_6 : std_logic_vector(1 downto 0);
  signal c_7 : std_logic_vector(1 downto 0);
  signal c_8 : std_logic_vector(1 downto 0);
  signal c_9 : std_logic_vector(1 downto 0);
  signal c_10 : std_logic_vector(1 downto 0);
  signal c_11 : std_logic_vector(1 downto 0);
  signal c_12 : std_logic_vector(1 downto 0);
  signal d_0 : std_logic_vector(1 downto 0);
  signal d_1 : std_logic_vector(1 downto 0);
  signal d_2 : std_logic_vector(1 downto 0);
  signal d_3 : std_logic_vector(1 downto 0);
  signal d_4 : std_logic_vector(1 downto 0);
  signal d_5 : std_logic_vector(1 downto 0);
  signal d_6 : std_logic_vector(1 downto 0);
  signal d_7 : std_logic_vector(1 downto 0);
  signal d_8 : std_logic_vector(1 downto 0);
  signal d_9 : std_logic_vector(1 downto 0);
  signal d_10 : std_logic_vector(1 downto 0);
  signal d_11 : std_logic_vector(1 downto 0);
  signal d_12 : std_logic_vector(1 downto 0);
  signal e_0 : std_logic_vector(1 downto 0);
  signal e_1 : std_logic_vector(1 downto 0);
  signal e_2 : std_logic_vector(1 downto 0);
  signal e_3 : std_logic_vector(1 downto 0);
  signal e_4 : std_logic_vector(1 downto 0);
  signal e_5 : std_logic_vector(1 downto 0);
  signal e_6 : std_logic_vector(1 downto 0);
  signal e_7 : std_logic_vector(1 downto 0);
  signal e_8 : std_logic_vector(1 downto 0);
  signal e_9 : std_logic_vector(1 downto 0);
  signal e_10 : std_logic_vector(1 downto 0);
  signal e_11 : std_logic_vector(1 downto 0);
  signal e_12 : std_logic_vector(1 downto 0);
  signal f_0 : std_logic_vector(1 downto 0);
  signal f_1 : std_logic_vector(1 downto 0);
  signal f_2 : std_logic_vector(1 downto 0);
  signal f_3 : std_logic_vector(1 downto 0);
  signal f_4 : std_logic_vector(1 downto 0);
  signal f_5 : std_logic_vector(1 downto 0);
  signal f_6 : std_logic_vector(1 downto 0);
  signal f_7 : std_logic_vector(1 downto 0);
  signal f_8 : std_logic_vector(1 downto 0);
  signal f_9 : std_logic_vector(1 downto 0);
  signal f_10 : std_logic_vector(1 downto 0);
  signal f_11 : std_logic_vector(1 downto 0);
  signal f_12 : std_logic_vector(1 downto 0);
  signal p_0 : std_logic_vector(1 downto 0);
  signal p_1 : std_logic_vector(1 downto 0);
  signal p_2 : std_logic_vector(1 downto 0);
  signal p_3 : std_logic_vector(1 downto 0);
  signal p_4 : std_logic_vector(1 downto 0);
  signal p_5 : std_logic_vector(1 downto 0);
  signal p_6 : std_logic_vector(1 downto 0);
  signal p_7 : std_logic_vector(1 downto 0);
  signal p_8 : std_logic_vector(1 downto 0);
  signal p_9 : std_logic_vector(1 downto 0);
  signal p_10 : std_logic_vector(1 downto 0);
  signal p_11 : std_logic_vector(1 downto 0);
  signal p_12 : std_logic_vector(1 downto 0);
  signal q_0 : std_logic_vector(1 downto 0);
  signal q_1 : std_logic_vector(1 downto 0);
  signal q_2 : std_logic_vector(1 downto 0);
  signal q_3 : std_logic_vector(1 downto 0);
  signal q_4 : std_logic_vector(1 downto 0);
  signal q_5 : std_logic_vector(1 downto 0);
  signal q_6 : std_logic_vector(1 downto 0);
  signal q_7 : std_logic_vector(1 downto 0);
  signal q_8 : std_logic_vector(1 downto 0);
  signal q_9 : std_logic_vector(1 downto 0);
  signal q_10 : std_logic_vector(1 downto 0);
  signal q_11 : std_logic_vector(1 downto 0);
  signal q_12 : std_logic_vector(1 downto 0);
begin
  mul1 : entity work.G4MulTIMaskedN
    port map ( 
      io_x_0 => a_0,
      io_x_1 => a_1,
      io_x_2 => a_2,
      io_x_3 => a_3,
      io_x_4 => a_4,
      io_x_5 => a_5,
      io_x_6 => a_6,
      io_x_7 => a_7,
      io_x_8 => a_8,
      io_x_9 => a_9,
      io_x_10 => a_10,
      io_x_11 => a_11,
      io_x_12 => a_12,
      io_y_0 => b_0,
      io_y_1 => b_1,
      io_y_2 => b_2,
      io_y_3 => b_3,
      io_y_4 => b_4,
      io_y_5 => b_5,
      io_y_6 => b_6,
      io_y_7 => b_7,
      io_y_8 => b_8,
      io_y_9 => b_9,
      io_y_10 => b_10,
      io_y_11 => b_11,
      io_y_12 => b_12,
      io_z_0 => mul1_io_z_0,
      io_z_1 => mul1_io_z_1,
      io_z_2 => mul1_io_z_2,
      io_z_3 => mul1_io_z_3,
      io_z_4 => mul1_io_z_4,
      io_z_5 => mul1_io_z_5,
      io_z_6 => mul1_io_z_6,
      io_z_7 => mul1_io_z_7,
      io_z_8 => mul1_io_z_8,
      io_z_9 => mul1_io_z_9,
      io_z_10 => mul1_io_z_10,
      io_z_11 => mul1_io_z_11,
      io_z_12 => mul1_io_z_12,
      clk => clk,
      reset => reset 
    );
  mul2 : entity work.G4MulTIMaskedN
    port map ( 
      io_x_0 => e_0,
      io_x_1 => e_1,
      io_x_2 => e_2,
      io_x_3 => e_3,
      io_x_4 => e_4,
      io_x_5 => e_5,
      io_x_6 => e_6,
      io_x_7 => e_7,
      io_x_8 => e_8,
      io_x_9 => e_9,
      io_x_10 => e_10,
      io_x_11 => e_11,
      io_x_12 => e_12,
      io_y_0 => b_0,
      io_y_1 => b_1,
      io_y_2 => b_2,
      io_y_3 => b_3,
      io_y_4 => b_4,
      io_y_5 => b_5,
      io_y_6 => b_6,
      io_y_7 => b_7,
      io_y_8 => b_8,
      io_y_9 => b_9,
      io_y_10 => b_10,
      io_y_11 => b_11,
      io_y_12 => b_12,
      io_z_0 => mul2_io_z_0,
      io_z_1 => mul2_io_z_1,
      io_z_2 => mul2_io_z_2,
      io_z_3 => mul2_io_z_3,
      io_z_4 => mul2_io_z_4,
      io_z_5 => mul2_io_z_5,
      io_z_6 => mul2_io_z_6,
      io_z_7 => mul2_io_z_7,
      io_z_8 => mul2_io_z_8,
      io_z_9 => mul2_io_z_9,
      io_z_10 => mul2_io_z_10,
      io_z_11 => mul2_io_z_11,
      io_z_12 => mul2_io_z_12,
      clk => clk,
      reset => reset 
    );
  mul3 : entity work.G4MulTIMaskedN
    port map ( 
      io_x_0 => e_0,
      io_x_1 => e_1,
      io_x_2 => e_2,
      io_x_3 => e_3,
      io_x_4 => e_4,
      io_x_5 => e_5,
      io_x_6 => e_6,
      io_x_7 => e_7,
      io_x_8 => e_8,
      io_x_9 => e_9,
      io_x_10 => e_10,
      io_x_11 => e_11,
      io_x_12 => e_12,
      io_y_0 => a_0,
      io_y_1 => a_1,
      io_y_2 => a_2,
      io_y_3 => a_3,
      io_y_4 => a_4,
      io_y_5 => a_5,
      io_y_6 => a_6,
      io_y_7 => a_7,
      io_y_8 => a_8,
      io_y_9 => a_9,
      io_y_10 => a_10,
      io_y_11 => a_11,
      io_y_12 => a_12,
      io_z_0 => mul3_io_z_0,
      io_z_1 => mul3_io_z_1,
      io_z_2 => mul3_io_z_2,
      io_z_3 => mul3_io_z_3,
      io_z_4 => mul3_io_z_4,
      io_z_5 => mul3_io_z_5,
      io_z_6 => mul3_io_z_6,
      io_z_7 => mul3_io_z_7,
      io_z_8 => mul3_io_z_8,
      io_z_9 => mul3_io_z_9,
      io_z_10 => mul3_io_z_10,
      io_z_11 => mul3_io_z_11,
      io_z_12 => mul3_io_z_12,
      clk => clk,
      reset => reset 
    );
  g4Sq_52 : entity work.G4Sq
    port map ( 
      io_t => f_0,
      io_x => g4Sq_52_io_x 
    );
  g4ScaleN_52 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_52_io_x,
      io_x => g4ScaleN_52_io_x 
    );
  g4Sq_53 : entity work.G4Sq
    port map ( 
      io_t => f_1,
      io_x => g4Sq_53_io_x 
    );
  g4ScaleN_53 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_53_io_x,
      io_x => g4ScaleN_53_io_x 
    );
  g4Sq_54 : entity work.G4Sq
    port map ( 
      io_t => f_2,
      io_x => g4Sq_54_io_x 
    );
  g4ScaleN_54 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_54_io_x,
      io_x => g4ScaleN_54_io_x 
    );
  g4Sq_55 : entity work.G4Sq
    port map ( 
      io_t => f_3,
      io_x => g4Sq_55_io_x 
    );
  g4ScaleN_55 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_55_io_x,
      io_x => g4ScaleN_55_io_x 
    );
  g4Sq_56 : entity work.G4Sq
    port map ( 
      io_t => f_4,
      io_x => g4Sq_56_io_x 
    );
  g4ScaleN_56 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_56_io_x,
      io_x => g4ScaleN_56_io_x 
    );
  g4Sq_57 : entity work.G4Sq
    port map ( 
      io_t => f_5,
      io_x => g4Sq_57_io_x 
    );
  g4ScaleN_57 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_57_io_x,
      io_x => g4ScaleN_57_io_x 
    );
  g4Sq_58 : entity work.G4Sq
    port map ( 
      io_t => f_6,
      io_x => g4Sq_58_io_x 
    );
  g4ScaleN_58 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_58_io_x,
      io_x => g4ScaleN_58_io_x 
    );
  g4Sq_59 : entity work.G4Sq
    port map ( 
      io_t => f_7,
      io_x => g4Sq_59_io_x 
    );
  g4ScaleN_59 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_59_io_x,
      io_x => g4ScaleN_59_io_x 
    );
  g4Sq_60 : entity work.G4Sq
    port map ( 
      io_t => f_8,
      io_x => g4Sq_60_io_x 
    );
  g4ScaleN_60 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_60_io_x,
      io_x => g4ScaleN_60_io_x 
    );
  g4Sq_61 : entity work.G4Sq
    port map ( 
      io_t => f_9,
      io_x => g4Sq_61_io_x 
    );
  g4ScaleN_61 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_61_io_x,
      io_x => g4ScaleN_61_io_x 
    );
  g4Sq_62 : entity work.G4Sq
    port map ( 
      io_t => f_10,
      io_x => g4Sq_62_io_x 
    );
  g4ScaleN_62 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_62_io_x,
      io_x => g4ScaleN_62_io_x 
    );
  g4Sq_63 : entity work.G4Sq
    port map ( 
      io_t => f_11,
      io_x => g4Sq_63_io_x 
    );
  g4ScaleN_63 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_63_io_x,
      io_x => g4ScaleN_63_io_x 
    );
  g4Sq_64 : entity work.G4Sq
    port map ( 
      io_t => f_12,
      io_x => g4Sq_64_io_x 
    );
  g4ScaleN_64 : entity work.G4ScaleN
    port map ( 
      io_t => g4Sq_64_io_x,
      io_x => g4ScaleN_64_io_x 
    );
  g4Sq_65 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_65_io_t,
      io_x => g4Sq_65_io_x 
    );
  g4Sq_66 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_66_io_t,
      io_x => g4Sq_66_io_x 
    );
  g4Sq_67 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_67_io_t,
      io_x => g4Sq_67_io_x 
    );
  g4Sq_68 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_68_io_t,
      io_x => g4Sq_68_io_x 
    );
  g4Sq_69 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_69_io_t,
      io_x => g4Sq_69_io_x 
    );
  g4Sq_70 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_70_io_t,
      io_x => g4Sq_70_io_x 
    );
  g4Sq_71 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_71_io_t,
      io_x => g4Sq_71_io_x 
    );
  g4Sq_72 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_72_io_t,
      io_x => g4Sq_72_io_x 
    );
  g4Sq_73 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_73_io_t,
      io_x => g4Sq_73_io_x 
    );
  g4Sq_74 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_74_io_t,
      io_x => g4Sq_74_io_x 
    );
  g4Sq_75 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_75_io_t,
      io_x => g4Sq_75_io_x 
    );
  g4Sq_76 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_76_io_t,
      io_x => g4Sq_76_io_x 
    );
  g4Sq_77 : entity work.G4Sq
    port map ( 
      io_t => g4Sq_77_io_t,
      io_x => g4Sq_77_io_x 
    );
  dummy <= pkg_toStdLogic(false);
  a_0 <= pkg_extract(io_x_0,3,2);
  b_0 <= pkg_extract(io_x_0,1,0);
  a_1 <= pkg_extract(io_x_1,3,2);
  b_1 <= pkg_extract(io_x_1,1,0);
  a_2 <= pkg_extract(io_x_2,3,2);
  b_2 <= pkg_extract(io_x_2,1,0);
  a_3 <= pkg_extract(io_x_3,3,2);
  b_3 <= pkg_extract(io_x_3,1,0);
  a_4 <= pkg_extract(io_x_4,3,2);
  b_4 <= pkg_extract(io_x_4,1,0);
  a_5 <= pkg_extract(io_x_5,3,2);
  b_5 <= pkg_extract(io_x_5,1,0);
  a_6 <= pkg_extract(io_x_6,3,2);
  b_6 <= pkg_extract(io_x_6,1,0);
  a_7 <= pkg_extract(io_x_7,3,2);
  b_7 <= pkg_extract(io_x_7,1,0);
  a_8 <= pkg_extract(io_x_8,3,2);
  b_8 <= pkg_extract(io_x_8,1,0);
  a_9 <= pkg_extract(io_x_9,3,2);
  b_9 <= pkg_extract(io_x_9,1,0);
  a_10 <= pkg_extract(io_x_10,3,2);
  b_10 <= pkg_extract(io_x_10,1,0);
  a_11 <= pkg_extract(io_x_11,3,2);
  b_11 <= pkg_extract(io_x_11,1,0);
  a_12 <= pkg_extract(io_x_12,3,2);
  b_12 <= pkg_extract(io_x_12,1,0);
  f_0 <= (a_0 xor b_0);
  f_1 <= (a_1 xor b_1);
  f_2 <= (a_2 xor b_2);
  f_3 <= (a_3 xor b_3);
  f_4 <= (a_4 xor b_4);
  f_5 <= (a_5 xor b_5);
  f_6 <= (a_6 xor b_6);
  f_7 <= (a_7 xor b_7);
  f_8 <= (a_8 xor b_8);
  f_9 <= (a_9 xor b_9);
  f_10 <= (a_10 xor b_10);
  f_11 <= (a_11 xor b_11);
  f_12 <= (a_12 xor b_12);
  d_0 <= mul1_io_z_0;
  d_1 <= mul1_io_z_1;
  d_2 <= mul1_io_z_2;
  d_3 <= mul1_io_z_3;
  d_4 <= mul1_io_z_4;
  d_5 <= mul1_io_z_5;
  d_6 <= mul1_io_z_6;
  d_7 <= mul1_io_z_7;
  d_8 <= mul1_io_z_8;
  d_9 <= mul1_io_z_9;
  d_10 <= mul1_io_z_10;
  d_11 <= mul1_io_z_11;
  d_12 <= mul1_io_z_12;
  c_0 <= g4ScaleN_52_io_x;
  c_1 <= g4ScaleN_53_io_x;
  c_2 <= g4ScaleN_54_io_x;
  c_3 <= g4ScaleN_55_io_x;
  c_4 <= g4ScaleN_56_io_x;
  c_5 <= g4ScaleN_57_io_x;
  c_6 <= g4ScaleN_58_io_x;
  c_7 <= g4ScaleN_59_io_x;
  c_8 <= g4ScaleN_60_io_x;
  c_9 <= g4ScaleN_61_io_x;
  c_10 <= g4ScaleN_62_io_x;
  c_11 <= g4ScaleN_63_io_x;
  c_12 <= g4ScaleN_64_io_x;
  g4Sq_65_io_t <= (c_0 xor d_0);
  e_0 <= g4Sq_65_io_x;
  g4Sq_66_io_t <= (c_1 xor d_1);
  e_1 <= g4Sq_66_io_x;
  g4Sq_67_io_t <= (c_2 xor d_2);
  e_2 <= g4Sq_67_io_x;
  g4Sq_68_io_t <= (c_3 xor d_3);
  e_3 <= g4Sq_68_io_x;
  g4Sq_69_io_t <= (c_4 xor d_4);
  e_4 <= g4Sq_69_io_x;
  g4Sq_70_io_t <= (c_5 xor d_5);
  e_5 <= g4Sq_70_io_x;
  g4Sq_71_io_t <= (c_6 xor d_6);
  e_6 <= g4Sq_71_io_x;
  g4Sq_72_io_t <= (c_7 xor d_7);
  e_7 <= g4Sq_72_io_x;
  g4Sq_73_io_t <= (c_8 xor d_8);
  e_8 <= g4Sq_73_io_x;
  g4Sq_74_io_t <= (c_9 xor d_9);
  e_9 <= g4Sq_74_io_x;
  g4Sq_75_io_t <= (c_10 xor d_10);
  e_10 <= g4Sq_75_io_x;
  g4Sq_76_io_t <= (c_11 xor d_11);
  e_11 <= g4Sq_76_io_x;
  g4Sq_77_io_t <= (c_12 xor d_12);
  e_12 <= g4Sq_77_io_x;
  p_0 <= mul2_io_z_0;
  p_1 <= mul2_io_z_1;
  p_2 <= mul2_io_z_2;
  p_3 <= mul2_io_z_3;
  p_4 <= mul2_io_z_4;
  p_5 <= mul2_io_z_5;
  p_6 <= mul2_io_z_6;
  p_7 <= mul2_io_z_7;
  p_8 <= mul2_io_z_8;
  p_9 <= mul2_io_z_9;
  p_10 <= mul2_io_z_10;
  p_11 <= mul2_io_z_11;
  p_12 <= mul2_io_z_12;
  q_0 <= mul3_io_z_0;
  q_1 <= mul3_io_z_1;
  q_2 <= mul3_io_z_2;
  q_3 <= mul3_io_z_3;
  q_4 <= mul3_io_z_4;
  q_5 <= mul3_io_z_5;
  q_6 <= mul3_io_z_6;
  q_7 <= mul3_io_z_7;
  q_8 <= mul3_io_z_8;
  q_9 <= mul3_io_z_9;
  q_10 <= mul3_io_z_10;
  q_11 <= mul3_io_z_11;
  q_12 <= mul3_io_z_12;
  io_z_0 <= pkg_cat(p_0,q_0);
  io_z_1 <= pkg_cat(p_1,q_1);
  io_z_2 <= pkg_cat(p_2,q_2);
  io_z_3 <= pkg_cat(p_3,q_3);
  io_z_4 <= pkg_cat(p_4,q_4);
  io_z_5 <= pkg_cat(p_5,q_5);
  io_z_6 <= pkg_cat(p_6,q_6);
  io_z_7 <= pkg_cat(p_7,q_7);
  io_z_8 <= pkg_cat(p_8,q_8);
  io_z_9 <= pkg_cat(p_9,q_9);
  io_z_10 <= pkg_cat(p_10,q_10);
  io_z_11 <= pkg_cat(p_11,q_11);
  io_z_12 <= pkg_cat(p_12,q_12);
end arch;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity G16SqSc is
  port(
    io_t : in std_logic_vector(3 downto 0);
    io_x : out std_logic_vector(3 downto 0)
  );
end G16SqSc;

architecture arch of G16SqSc is
  signal square1_io_t : std_logic_vector(1 downto 0);
  signal square1_io_x : std_logic_vector(1 downto 0);
  signal square2_io_x : std_logic_vector(1 downto 0);
  signal scale_io_x : std_logic_vector(1 downto 0);

  signal a : std_logic_vector(1 downto 0);
  signal b : std_logic_vector(1 downto 0);
  signal c : std_logic_vector(1 downto 0);
  signal p : std_logic_vector(1 downto 0);
  signal q : std_logic_vector(1 downto 0);
begin
  square1 : entity work.G4Sq
    port map ( 
      io_t => square1_io_t,
      io_x => square1_io_x 
    );
  square2 : entity work.G4Sq
    port map ( 
      io_t => b,
      io_x => square2_io_x 
    );
  scale : entity work.G4ScaleN2
    port map ( 
      io_t => c,
      io_x => scale_io_x 
    );
  square1_io_t <= (a xor b);
  p <= square1_io_x;
  c <= square2_io_x;
  q <= scale_io_x;
  a <= pkg_extract(io_t,3,2);
  b <= pkg_extract(io_t,1,0);
  io_x <= pkg_cat(p,q);
end arch;


--G16SqSc_1 replaced by G16SqSc


--G16SqSc_2 replaced by G16SqSc


--G16SqSc_3 replaced by G16SqSc


--G16SqSc_4 replaced by G16SqSc


--G16SqSc_5 replaced by G16SqSc


--G16SqSc_6 replaced by G16SqSc


--G16SqSc_7 replaced by G16SqSc


--G16SqSc_8 replaced by G16SqSc


--G16SqSc_9 replaced by G16SqSc


--G16SqSc_10 replaced by G16SqSc


--G16SqSc_11 replaced by G16SqSc


--G16SqSc_12 replaced by G16SqSc

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg_scala2hdl.all;
use work.all;
use work.pkg_enum.all;


entity G256InvTIMaskedN is
  port(
    io_x_0 : in std_logic_vector(7 downto 0);
    io_x_1 : in std_logic_vector(7 downto 0);
    io_x_2 : in std_logic_vector(7 downto 0);
    io_x_3 : in std_logic_vector(7 downto 0);
    io_x_4 : in std_logic_vector(7 downto 0);
    io_x_5 : in std_logic_vector(7 downto 0);
    io_x_6 : in std_logic_vector(7 downto 0);
    io_x_7 : in std_logic_vector(7 downto 0);
    io_x_8 : in std_logic_vector(7 downto 0);
    io_x_9 : in std_logic_vector(7 downto 0);
    io_x_10 : in std_logic_vector(7 downto 0);
    io_x_11 : in std_logic_vector(7 downto 0);
    io_x_12 : in std_logic_vector(7 downto 0);
    io_z_0 : out std_logic_vector(7 downto 0);
    io_z_1 : out std_logic_vector(7 downto 0);
    io_z_2 : out std_logic_vector(7 downto 0);
    io_z_3 : out std_logic_vector(7 downto 0);
    io_z_4 : out std_logic_vector(7 downto 0);
    io_z_5 : out std_logic_vector(7 downto 0);
    io_z_6 : out std_logic_vector(7 downto 0);
    io_z_7 : out std_logic_vector(7 downto 0);
    io_z_8 : out std_logic_vector(7 downto 0);
    io_z_9 : out std_logic_vector(7 downto 0);
    io_z_10 : out std_logic_vector(7 downto 0);
    io_z_11 : out std_logic_vector(7 downto 0);
    io_z_12 : out std_logic_vector(7 downto 0);
    clk : in std_logic;
    reset : in std_logic
  );
end G256InvTIMaskedN;

architecture arch of G256InvTIMaskedN is
  signal inv_io_x_0 : std_logic_vector(3 downto 0);
  signal inv_io_x_1 : std_logic_vector(3 downto 0);
  signal inv_io_x_2 : std_logic_vector(3 downto 0);
  signal inv_io_x_3 : std_logic_vector(3 downto 0);
  signal inv_io_x_4 : std_logic_vector(3 downto 0);
  signal inv_io_x_5 : std_logic_vector(3 downto 0);
  signal inv_io_x_6 : std_logic_vector(3 downto 0);
  signal inv_io_x_7 : std_logic_vector(3 downto 0);
  signal inv_io_x_8 : std_logic_vector(3 downto 0);
  signal inv_io_x_9 : std_logic_vector(3 downto 0);
  signal inv_io_x_10 : std_logic_vector(3 downto 0);
  signal inv_io_x_11 : std_logic_vector(3 downto 0);
  signal inv_io_x_12 : std_logic_vector(3 downto 0);
  signal mul1_io_z_0 : std_logic_vector(3 downto 0);
  signal mul1_io_z_1 : std_logic_vector(3 downto 0);
  signal mul1_io_z_2 : std_logic_vector(3 downto 0);
  signal mul1_io_z_3 : std_logic_vector(3 downto 0);
  signal mul1_io_z_4 : std_logic_vector(3 downto 0);
  signal mul1_io_z_5 : std_logic_vector(3 downto 0);
  signal mul1_io_z_6 : std_logic_vector(3 downto 0);
  signal mul1_io_z_7 : std_logic_vector(3 downto 0);
  signal mul1_io_z_8 : std_logic_vector(3 downto 0);
  signal mul1_io_z_9 : std_logic_vector(3 downto 0);
  signal mul1_io_z_10 : std_logic_vector(3 downto 0);
  signal mul1_io_z_11 : std_logic_vector(3 downto 0);
  signal mul1_io_z_12 : std_logic_vector(3 downto 0);
  signal mul2_io_z_0 : std_logic_vector(3 downto 0);
  signal mul2_io_z_1 : std_logic_vector(3 downto 0);
  signal mul2_io_z_2 : std_logic_vector(3 downto 0);
  signal mul2_io_z_3 : std_logic_vector(3 downto 0);
  signal mul2_io_z_4 : std_logic_vector(3 downto 0);
  signal mul2_io_z_5 : std_logic_vector(3 downto 0);
  signal mul2_io_z_6 : std_logic_vector(3 downto 0);
  signal mul2_io_z_7 : std_logic_vector(3 downto 0);
  signal mul2_io_z_8 : std_logic_vector(3 downto 0);
  signal mul2_io_z_9 : std_logic_vector(3 downto 0);
  signal mul2_io_z_10 : std_logic_vector(3 downto 0);
  signal mul2_io_z_11 : std_logic_vector(3 downto 0);
  signal mul2_io_z_12 : std_logic_vector(3 downto 0);
  signal mul3_io_z_0 : std_logic_vector(3 downto 0);
  signal mul3_io_z_1 : std_logic_vector(3 downto 0);
  signal mul3_io_z_2 : std_logic_vector(3 downto 0);
  signal mul3_io_z_3 : std_logic_vector(3 downto 0);
  signal mul3_io_z_4 : std_logic_vector(3 downto 0);
  signal mul3_io_z_5 : std_logic_vector(3 downto 0);
  signal mul3_io_z_6 : std_logic_vector(3 downto 0);
  signal mul3_io_z_7 : std_logic_vector(3 downto 0);
  signal mul3_io_z_8 : std_logic_vector(3 downto 0);
  signal mul3_io_z_9 : std_logic_vector(3 downto 0);
  signal mul3_io_z_10 : std_logic_vector(3 downto 0);
  signal mul3_io_z_11 : std_logic_vector(3 downto 0);
  signal mul3_io_z_12 : std_logic_vector(3 downto 0);
  signal inv_io_z_0 : std_logic_vector(3 downto 0);
  signal inv_io_z_1 : std_logic_vector(3 downto 0);
  signal inv_io_z_2 : std_logic_vector(3 downto 0);
  signal inv_io_z_3 : std_logic_vector(3 downto 0);
  signal inv_io_z_4 : std_logic_vector(3 downto 0);
  signal inv_io_z_5 : std_logic_vector(3 downto 0);
  signal inv_io_z_6 : std_logic_vector(3 downto 0);
  signal inv_io_z_7 : std_logic_vector(3 downto 0);
  signal inv_io_z_8 : std_logic_vector(3 downto 0);
  signal inv_io_z_9 : std_logic_vector(3 downto 0);
  signal inv_io_z_10 : std_logic_vector(3 downto 0);
  signal inv_io_z_11 : std_logic_vector(3 downto 0);
  signal inv_io_z_12 : std_logic_vector(3 downto 0);
  signal g16SqSc_13_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_14_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_15_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_16_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_17_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_18_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_19_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_20_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_21_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_22_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_23_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_24_io_x : std_logic_vector(3 downto 0);
  signal g16SqSc_25_io_x : std_logic_vector(3 downto 0);

  signal dummy : std_logic;
  signal a_0 : std_logic_vector(3 downto 0);
  signal a_1 : std_logic_vector(3 downto 0);
  signal a_2 : std_logic_vector(3 downto 0);
  signal a_3 : std_logic_vector(3 downto 0);
  signal a_4 : std_logic_vector(3 downto 0);
  signal a_5 : std_logic_vector(3 downto 0);
  signal a_6 : std_logic_vector(3 downto 0);
  signal a_7 : std_logic_vector(3 downto 0);
  signal a_8 : std_logic_vector(3 downto 0);
  signal a_9 : std_logic_vector(3 downto 0);
  signal a_10 : std_logic_vector(3 downto 0);
  signal a_11 : std_logic_vector(3 downto 0);
  signal a_12 : std_logic_vector(3 downto 0);
  signal b_0 : std_logic_vector(3 downto 0);
  signal b_1 : std_logic_vector(3 downto 0);
  signal b_2 : std_logic_vector(3 downto 0);
  signal b_3 : std_logic_vector(3 downto 0);
  signal b_4 : std_logic_vector(3 downto 0);
  signal b_5 : std_logic_vector(3 downto 0);
  signal b_6 : std_logic_vector(3 downto 0);
  signal b_7 : std_logic_vector(3 downto 0);
  signal b_8 : std_logic_vector(3 downto 0);
  signal b_9 : std_logic_vector(3 downto 0);
  signal b_10 : std_logic_vector(3 downto 0);
  signal b_11 : std_logic_vector(3 downto 0);
  signal b_12 : std_logic_vector(3 downto 0);
  signal c_0 : std_logic_vector(3 downto 0);
  signal c_1 : std_logic_vector(3 downto 0);
  signal c_2 : std_logic_vector(3 downto 0);
  signal c_3 : std_logic_vector(3 downto 0);
  signal c_4 : std_logic_vector(3 downto 0);
  signal c_5 : std_logic_vector(3 downto 0);
  signal c_6 : std_logic_vector(3 downto 0);
  signal c_7 : std_logic_vector(3 downto 0);
  signal c_8 : std_logic_vector(3 downto 0);
  signal c_9 : std_logic_vector(3 downto 0);
  signal c_10 : std_logic_vector(3 downto 0);
  signal c_11 : std_logic_vector(3 downto 0);
  signal c_12 : std_logic_vector(3 downto 0);
  signal d_0 : std_logic_vector(3 downto 0);
  signal d_1 : std_logic_vector(3 downto 0);
  signal d_2 : std_logic_vector(3 downto 0);
  signal d_3 : std_logic_vector(3 downto 0);
  signal d_4 : std_logic_vector(3 downto 0);
  signal d_5 : std_logic_vector(3 downto 0);
  signal d_6 : std_logic_vector(3 downto 0);
  signal d_7 : std_logic_vector(3 downto 0);
  signal d_8 : std_logic_vector(3 downto 0);
  signal d_9 : std_logic_vector(3 downto 0);
  signal d_10 : std_logic_vector(3 downto 0);
  signal d_11 : std_logic_vector(3 downto 0);
  signal d_12 : std_logic_vector(3 downto 0);
  signal e_0 : std_logic_vector(3 downto 0);
  signal e_1 : std_logic_vector(3 downto 0);
  signal e_2 : std_logic_vector(3 downto 0);
  signal e_3 : std_logic_vector(3 downto 0);
  signal e_4 : std_logic_vector(3 downto 0);
  signal e_5 : std_logic_vector(3 downto 0);
  signal e_6 : std_logic_vector(3 downto 0);
  signal e_7 : std_logic_vector(3 downto 0);
  signal e_8 : std_logic_vector(3 downto 0);
  signal e_9 : std_logic_vector(3 downto 0);
  signal e_10 : std_logic_vector(3 downto 0);
  signal e_11 : std_logic_vector(3 downto 0);
  signal e_12 : std_logic_vector(3 downto 0);
  signal f_0 : std_logic_vector(3 downto 0);
  signal f_1 : std_logic_vector(3 downto 0);
  signal f_2 : std_logic_vector(3 downto 0);
  signal f_3 : std_logic_vector(3 downto 0);
  signal f_4 : std_logic_vector(3 downto 0);
  signal f_5 : std_logic_vector(3 downto 0);
  signal f_6 : std_logic_vector(3 downto 0);
  signal f_7 : std_logic_vector(3 downto 0);
  signal f_8 : std_logic_vector(3 downto 0);
  signal f_9 : std_logic_vector(3 downto 0);
  signal f_10 : std_logic_vector(3 downto 0);
  signal f_11 : std_logic_vector(3 downto 0);
  signal f_12 : std_logic_vector(3 downto 0);
  signal p_0 : std_logic_vector(3 downto 0);
  signal p_1 : std_logic_vector(3 downto 0);
  signal p_2 : std_logic_vector(3 downto 0);
  signal p_3 : std_logic_vector(3 downto 0);
  signal p_4 : std_logic_vector(3 downto 0);
  signal p_5 : std_logic_vector(3 downto 0);
  signal p_6 : std_logic_vector(3 downto 0);
  signal p_7 : std_logic_vector(3 downto 0);
  signal p_8 : std_logic_vector(3 downto 0);
  signal p_9 : std_logic_vector(3 downto 0);
  signal p_10 : std_logic_vector(3 downto 0);
  signal p_11 : std_logic_vector(3 downto 0);
  signal p_12 : std_logic_vector(3 downto 0);
  signal q_0 : std_logic_vector(3 downto 0);
  signal q_1 : std_logic_vector(3 downto 0);
  signal q_2 : std_logic_vector(3 downto 0);
  signal q_3 : std_logic_vector(3 downto 0);
  signal q_4 : std_logic_vector(3 downto 0);
  signal q_5 : std_logic_vector(3 downto 0);
  signal q_6 : std_logic_vector(3 downto 0);
  signal q_7 : std_logic_vector(3 downto 0);
  signal q_8 : std_logic_vector(3 downto 0);
  signal q_9 : std_logic_vector(3 downto 0);
  signal q_10 : std_logic_vector(3 downto 0);
  signal q_11 : std_logic_vector(3 downto 0);
  signal q_12 : std_logic_vector(3 downto 0);
begin
  mul1 : entity work.G16MulTIMaskedN
    port map ( 
      io_x_0 => a_0,
      io_x_1 => a_1,
      io_x_2 => a_2,
      io_x_3 => a_3,
      io_x_4 => a_4,
      io_x_5 => a_5,
      io_x_6 => a_6,
      io_x_7 => a_7,
      io_x_8 => a_8,
      io_x_9 => a_9,
      io_x_10 => a_10,
      io_x_11 => a_11,
      io_x_12 => a_12,
      io_y_0 => b_0,
      io_y_1 => b_1,
      io_y_2 => b_2,
      io_y_3 => b_3,
      io_y_4 => b_4,
      io_y_5 => b_5,
      io_y_6 => b_6,
      io_y_7 => b_7,
      io_y_8 => b_8,
      io_y_9 => b_9,
      io_y_10 => b_10,
      io_y_11 => b_11,
      io_y_12 => b_12,
      io_z_0 => mul1_io_z_0,
      io_z_1 => mul1_io_z_1,
      io_z_2 => mul1_io_z_2,
      io_z_3 => mul1_io_z_3,
      io_z_4 => mul1_io_z_4,
      io_z_5 => mul1_io_z_5,
      io_z_6 => mul1_io_z_6,
      io_z_7 => mul1_io_z_7,
      io_z_8 => mul1_io_z_8,
      io_z_9 => mul1_io_z_9,
      io_z_10 => mul1_io_z_10,
      io_z_11 => mul1_io_z_11,
      io_z_12 => mul1_io_z_12,
      clk => clk,
      reset => reset 
    );
  mul2 : entity work.G16MulTIMaskedN
    port map ( 
      io_x_0 => e_0,
      io_x_1 => e_1,
      io_x_2 => e_2,
      io_x_3 => e_3,
      io_x_4 => e_4,
      io_x_5 => e_5,
      io_x_6 => e_6,
      io_x_7 => e_7,
      io_x_8 => e_8,
      io_x_9 => e_9,
      io_x_10 => e_10,
      io_x_11 => e_11,
      io_x_12 => e_12,
      io_y_0 => b_0,
      io_y_1 => b_1,
      io_y_2 => b_2,
      io_y_3 => b_3,
      io_y_4 => b_4,
      io_y_5 => b_5,
      io_y_6 => b_6,
      io_y_7 => b_7,
      io_y_8 => b_8,
      io_y_9 => b_9,
      io_y_10 => b_10,
      io_y_11 => b_11,
      io_y_12 => b_12,
      io_z_0 => mul2_io_z_0,
      io_z_1 => mul2_io_z_1,
      io_z_2 => mul2_io_z_2,
      io_z_3 => mul2_io_z_3,
      io_z_4 => mul2_io_z_4,
      io_z_5 => mul2_io_z_5,
      io_z_6 => mul2_io_z_6,
      io_z_7 => mul2_io_z_7,
      io_z_8 => mul2_io_z_8,
      io_z_9 => mul2_io_z_9,
      io_z_10 => mul2_io_z_10,
      io_z_11 => mul2_io_z_11,
      io_z_12 => mul2_io_z_12,
      clk => clk,
      reset => reset 
    );
  mul3 : entity work.G16MulTIMaskedN
    port map ( 
      io_x_0 => e_0,
      io_x_1 => e_1,
      io_x_2 => e_2,
      io_x_3 => e_3,
      io_x_4 => e_4,
      io_x_5 => e_5,
      io_x_6 => e_6,
      io_x_7 => e_7,
      io_x_8 => e_8,
      io_x_9 => e_9,
      io_x_10 => e_10,
      io_x_11 => e_11,
      io_x_12 => e_12,
      io_y_0 => a_0,
      io_y_1 => a_1,
      io_y_2 => a_2,
      io_y_3 => a_3,
      io_y_4 => a_4,
      io_y_5 => a_5,
      io_y_6 => a_6,
      io_y_7 => a_7,
      io_y_8 => a_8,
      io_y_9 => a_9,
      io_y_10 => a_10,
      io_y_11 => a_11,
      io_y_12 => a_12,
      io_z_0 => mul3_io_z_0,
      io_z_1 => mul3_io_z_1,
      io_z_2 => mul3_io_z_2,
      io_z_3 => mul3_io_z_3,
      io_z_4 => mul3_io_z_4,
      io_z_5 => mul3_io_z_5,
      io_z_6 => mul3_io_z_6,
      io_z_7 => mul3_io_z_7,
      io_z_8 => mul3_io_z_8,
      io_z_9 => mul3_io_z_9,
      io_z_10 => mul3_io_z_10,
      io_z_11 => mul3_io_z_11,
      io_z_12 => mul3_io_z_12,
      clk => clk,
      reset => reset 
    );
  inv : entity work.G16InvTIMaskedN
    port map ( 
      io_x_0 => inv_io_x_0,
      io_x_1 => inv_io_x_1,
      io_x_2 => inv_io_x_2,
      io_x_3 => inv_io_x_3,
      io_x_4 => inv_io_x_4,
      io_x_5 => inv_io_x_5,
      io_x_6 => inv_io_x_6,
      io_x_7 => inv_io_x_7,
      io_x_8 => inv_io_x_8,
      io_x_9 => inv_io_x_9,
      io_x_10 => inv_io_x_10,
      io_x_11 => inv_io_x_11,
      io_x_12 => inv_io_x_12,
      io_z_0 => inv_io_z_0,
      io_z_1 => inv_io_z_1,
      io_z_2 => inv_io_z_2,
      io_z_3 => inv_io_z_3,
      io_z_4 => inv_io_z_4,
      io_z_5 => inv_io_z_5,
      io_z_6 => inv_io_z_6,
      io_z_7 => inv_io_z_7,
      io_z_8 => inv_io_z_8,
      io_z_9 => inv_io_z_9,
      io_z_10 => inv_io_z_10,
      io_z_11 => inv_io_z_11,
      io_z_12 => inv_io_z_12,
      clk => clk,
      reset => reset 
    );
  g16SqSc_13 : entity work.G16SqSc
    port map ( 
      io_t => f_0,
      io_x => g16SqSc_13_io_x 
    );
  g16SqSc_14 : entity work.G16SqSc
    port map ( 
      io_t => f_1,
      io_x => g16SqSc_14_io_x 
    );
  g16SqSc_15 : entity work.G16SqSc
    port map ( 
      io_t => f_2,
      io_x => g16SqSc_15_io_x 
    );
  g16SqSc_16 : entity work.G16SqSc
    port map ( 
      io_t => f_3,
      io_x => g16SqSc_16_io_x 
    );
  g16SqSc_17 : entity work.G16SqSc
    port map ( 
      io_t => f_4,
      io_x => g16SqSc_17_io_x 
    );
  g16SqSc_18 : entity work.G16SqSc
    port map ( 
      io_t => f_5,
      io_x => g16SqSc_18_io_x 
    );
  g16SqSc_19 : entity work.G16SqSc
    port map ( 
      io_t => f_6,
      io_x => g16SqSc_19_io_x 
    );
  g16SqSc_20 : entity work.G16SqSc
    port map ( 
      io_t => f_7,
      io_x => g16SqSc_20_io_x 
    );
  g16SqSc_21 : entity work.G16SqSc
    port map ( 
      io_t => f_8,
      io_x => g16SqSc_21_io_x 
    );
  g16SqSc_22 : entity work.G16SqSc
    port map ( 
      io_t => f_9,
      io_x => g16SqSc_22_io_x 
    );
  g16SqSc_23 : entity work.G16SqSc
    port map ( 
      io_t => f_10,
      io_x => g16SqSc_23_io_x 
    );
  g16SqSc_24 : entity work.G16SqSc
    port map ( 
      io_t => f_11,
      io_x => g16SqSc_24_io_x 
    );
  g16SqSc_25 : entity work.G16SqSc
    port map ( 
      io_t => f_12,
      io_x => g16SqSc_25_io_x 
    );
  dummy <= pkg_toStdLogic(false);
  a_0 <= pkg_extract(io_x_0,7,4);
  b_0 <= pkg_extract(io_x_0,3,0);
  a_1 <= pkg_extract(io_x_1,7,4);
  b_1 <= pkg_extract(io_x_1,3,0);
  a_2 <= pkg_extract(io_x_2,7,4);
  b_2 <= pkg_extract(io_x_2,3,0);
  a_3 <= pkg_extract(io_x_3,7,4);
  b_3 <= pkg_extract(io_x_3,3,0);
  a_4 <= pkg_extract(io_x_4,7,4);
  b_4 <= pkg_extract(io_x_4,3,0);
  a_5 <= pkg_extract(io_x_5,7,4);
  b_5 <= pkg_extract(io_x_5,3,0);
  a_6 <= pkg_extract(io_x_6,7,4);
  b_6 <= pkg_extract(io_x_6,3,0);
  a_7 <= pkg_extract(io_x_7,7,4);
  b_7 <= pkg_extract(io_x_7,3,0);
  a_8 <= pkg_extract(io_x_8,7,4);
  b_8 <= pkg_extract(io_x_8,3,0);
  a_9 <= pkg_extract(io_x_9,7,4);
  b_9 <= pkg_extract(io_x_9,3,0);
  a_10 <= pkg_extract(io_x_10,7,4);
  b_10 <= pkg_extract(io_x_10,3,0);
  a_11 <= pkg_extract(io_x_11,7,4);
  b_11 <= pkg_extract(io_x_11,3,0);
  a_12 <= pkg_extract(io_x_12,7,4);
  b_12 <= pkg_extract(io_x_12,3,0);
  f_0 <= (a_0 xor b_0);
  f_1 <= (a_1 xor b_1);
  f_2 <= (a_2 xor b_2);
  f_3 <= (a_3 xor b_3);
  f_4 <= (a_4 xor b_4);
  f_5 <= (a_5 xor b_5);
  f_6 <= (a_6 xor b_6);
  f_7 <= (a_7 xor b_7);
  f_8 <= (a_8 xor b_8);
  f_9 <= (a_9 xor b_9);
  f_10 <= (a_10 xor b_10);
  f_11 <= (a_11 xor b_11);
  f_12 <= (a_12 xor b_12);
  c_0 <= g16SqSc_13_io_x;
  c_1 <= g16SqSc_14_io_x;
  c_2 <= g16SqSc_15_io_x;
  c_3 <= g16SqSc_16_io_x;
  c_4 <= g16SqSc_17_io_x;
  c_5 <= g16SqSc_18_io_x;
  c_6 <= g16SqSc_19_io_x;
  c_7 <= g16SqSc_20_io_x;
  c_8 <= g16SqSc_21_io_x;
  c_9 <= g16SqSc_22_io_x;
  c_10 <= g16SqSc_23_io_x;
  c_11 <= g16SqSc_24_io_x;
  c_12 <= g16SqSc_25_io_x;
  d_0 <= mul1_io_z_0;
  d_1 <= mul1_io_z_1;
  d_2 <= mul1_io_z_2;
  d_3 <= mul1_io_z_3;
  d_4 <= mul1_io_z_4;
  d_5 <= mul1_io_z_5;
  d_6 <= mul1_io_z_6;
  d_7 <= mul1_io_z_7;
  d_8 <= mul1_io_z_8;
  d_9 <= mul1_io_z_9;
  d_10 <= mul1_io_z_10;
  d_11 <= mul1_io_z_11;
  d_12 <= mul1_io_z_12;
  inv_io_x_0 <= (c_0 xor d_0);
  inv_io_x_1 <= (c_1 xor d_1);
  inv_io_x_2 <= (c_2 xor d_2);
  inv_io_x_3 <= (c_3 xor d_3);
  inv_io_x_4 <= (c_4 xor d_4);
  inv_io_x_5 <= (c_5 xor d_5);
  inv_io_x_6 <= (c_6 xor d_6);
  inv_io_x_7 <= (c_7 xor d_7);
  inv_io_x_8 <= (c_8 xor d_8);
  inv_io_x_9 <= (c_9 xor d_9);
  inv_io_x_10 <= (c_10 xor d_10);
  inv_io_x_11 <= (c_11 xor d_11);
  inv_io_x_12 <= (c_12 xor d_12);
  e_0 <= inv_io_z_0;
  e_1 <= inv_io_z_1;
  e_2 <= inv_io_z_2;
  e_3 <= inv_io_z_3;
  e_4 <= inv_io_z_4;
  e_5 <= inv_io_z_5;
  e_6 <= inv_io_z_6;
  e_7 <= inv_io_z_7;
  e_8 <= inv_io_z_8;
  e_9 <= inv_io_z_9;
  e_10 <= inv_io_z_10;
  e_11 <= inv_io_z_11;
  e_12 <= inv_io_z_12;
  p_0 <= mul2_io_z_0;
  p_1 <= mul2_io_z_1;
  p_2 <= mul2_io_z_2;
  p_3 <= mul2_io_z_3;
  p_4 <= mul2_io_z_4;
  p_5 <= mul2_io_z_5;
  p_6 <= mul2_io_z_6;
  p_7 <= mul2_io_z_7;
  p_8 <= mul2_io_z_8;
  p_9 <= mul2_io_z_9;
  p_10 <= mul2_io_z_10;
  p_11 <= mul2_io_z_11;
  p_12 <= mul2_io_z_12;
  q_0 <= mul3_io_z_0;
  q_1 <= mul3_io_z_1;
  q_2 <= mul3_io_z_2;
  q_3 <= mul3_io_z_3;
  q_4 <= mul3_io_z_4;
  q_5 <= mul3_io_z_5;
  q_6 <= mul3_io_z_6;
  q_7 <= mul3_io_z_7;
  q_8 <= mul3_io_z_8;
  q_9 <= mul3_io_z_9;
  q_10 <= mul3_io_z_10;
  q_11 <= mul3_io_z_11;
  q_12 <= mul3_io_z_12;
  io_z_0 <= pkg_cat(p_0,q_0);
  io_z_1 <= pkg_cat(p_1,q_1);
  io_z_2 <= pkg_cat(p_2,q_2);
  io_z_3 <= pkg_cat(p_3,q_3);
  io_z_4 <= pkg_cat(p_4,q_4);
  io_z_5 <= pkg_cat(p_5,q_5);
  io_z_6 <= pkg_cat(p_6,q_6);
  io_z_7 <= pkg_cat(p_7,q_7);
  io_z_8 <= pkg_cat(p_8,q_8);
  io_z_9 <= pkg_cat(p_9,q_9);
  io_z_10 <= pkg_cat(p_10,q_10);
  io_z_11 <= pkg_cat(p_11,q_11);
  io_z_12 <= pkg_cat(p_12,q_12);
end arch;

