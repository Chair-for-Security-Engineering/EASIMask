// Generator : SpinalHDL v1.6.2    git head : 685405804ac0fa51f884fe0ee6813ba6f1f31e4e
// Component : aesEncrypt
// Git hash  : 685405804ac0fa51f884fe0ee6813ba6f1f31e4e

`timescale 1ns/1ps 

module aesEncrypt (
  input               io_reset,
  input      [127:0]  io_pt,
  input      [127:0]  io_key,
  output reg [127:0]  io_ret,
  output reg          io_done,
  input               clk,
  input               reset
);
  localparam fsm_enumDef_BOOT = 2'd0;
  localparam fsm_enumDef_sReset = 2'd1;
  localparam fsm_enumDef_sAESRound = 2'd2;
  localparam fsm_enumDef_sAESFinalRound = 2'd3;

  reg        [7:0]    addroundkey_1_io_rk_0_0;
  reg        [7:0]    addroundkey_1_io_rk_0_1;
  reg        [7:0]    addroundkey_1_io_rk_0_2;
  reg        [7:0]    addroundkey_1_io_rk_0_3;
  reg        [7:0]    addroundkey_1_io_rk_1_0;
  reg        [7:0]    addroundkey_1_io_rk_1_1;
  reg        [7:0]    addroundkey_1_io_rk_1_2;
  reg        [7:0]    addroundkey_1_io_rk_1_3;
  reg        [7:0]    addroundkey_1_io_rk_2_0;
  reg        [7:0]    addroundkey_1_io_rk_2_1;
  reg        [7:0]    addroundkey_1_io_rk_2_2;
  reg        [7:0]    addroundkey_1_io_rk_2_3;
  reg        [7:0]    addroundkey_1_io_rk_3_0;
  reg        [7:0]    addroundkey_1_io_rk_3_1;
  reg        [7:0]    addroundkey_1_io_rk_3_2;
  reg        [7:0]    addroundkey_1_io_rk_3_3;
  reg        [7:0]    addroundkey_1_io_s_0_0;
  reg        [7:0]    addroundkey_1_io_s_0_1;
  reg        [7:0]    addroundkey_1_io_s_0_2;
  reg        [7:0]    addroundkey_1_io_s_0_3;
  reg        [7:0]    addroundkey_1_io_s_1_0;
  reg        [7:0]    addroundkey_1_io_s_1_1;
  reg        [7:0]    addroundkey_1_io_s_1_2;
  reg        [7:0]    addroundkey_1_io_s_1_3;
  reg        [7:0]    addroundkey_1_io_s_2_0;
  reg        [7:0]    addroundkey_1_io_s_2_1;
  reg        [7:0]    addroundkey_1_io_s_2_2;
  reg        [7:0]    addroundkey_1_io_s_2_3;
  reg        [7:0]    addroundkey_1_io_s_3_0;
  reg        [7:0]    addroundkey_1_io_s_3_1;
  reg        [7:0]    addroundkey_1_io_s_3_2;
  reg        [7:0]    addroundkey_1_io_s_3_3;
  reg        [7:0]    keyschedule_1_io_key_0_0;
  reg        [7:0]    keyschedule_1_io_key_0_1;
  reg        [7:0]    keyschedule_1_io_key_0_2;
  reg        [7:0]    keyschedule_1_io_key_0_3;
  reg        [7:0]    keyschedule_1_io_key_1_0;
  reg        [7:0]    keyschedule_1_io_key_1_1;
  reg        [7:0]    keyschedule_1_io_key_1_2;
  reg        [7:0]    keyschedule_1_io_key_1_3;
  reg        [7:0]    keyschedule_1_io_key_2_0;
  reg        [7:0]    keyschedule_1_io_key_2_1;
  reg        [7:0]    keyschedule_1_io_key_2_2;
  reg        [7:0]    keyschedule_1_io_key_2_3;
  reg        [7:0]    keyschedule_1_io_key_3_0;
  reg        [7:0]    keyschedule_1_io_key_3_1;
  reg        [7:0]    keyschedule_1_io_key_3_2;
  reg        [7:0]    keyschedule_1_io_key_3_3;
  wire       [7:0]    addroundkey_1_io_ret_0_0;
  wire       [7:0]    addroundkey_1_io_ret_0_1;
  wire       [7:0]    addroundkey_1_io_ret_0_2;
  wire       [7:0]    addroundkey_1_io_ret_0_3;
  wire       [7:0]    addroundkey_1_io_ret_1_0;
  wire       [7:0]    addroundkey_1_io_ret_1_1;
  wire       [7:0]    addroundkey_1_io_ret_1_2;
  wire       [7:0]    addroundkey_1_io_ret_1_3;
  wire       [7:0]    addroundkey_1_io_ret_2_0;
  wire       [7:0]    addroundkey_1_io_ret_2_1;
  wire       [7:0]    addroundkey_1_io_ret_2_2;
  wire       [7:0]    addroundkey_1_io_ret_2_3;
  wire       [7:0]    addroundkey_1_io_ret_3_0;
  wire       [7:0]    addroundkey_1_io_ret_3_1;
  wire       [7:0]    addroundkey_1_io_ret_3_2;
  wire       [7:0]    addroundkey_1_io_ret_3_3;
  wire       [7:0]    subbytes_1_io_ret_0_0;
  wire       [7:0]    subbytes_1_io_ret_0_1;
  wire       [7:0]    subbytes_1_io_ret_0_2;
  wire       [7:0]    subbytes_1_io_ret_0_3;
  wire       [7:0]    subbytes_1_io_ret_1_0;
  wire       [7:0]    subbytes_1_io_ret_1_1;
  wire       [7:0]    subbytes_1_io_ret_1_2;
  wire       [7:0]    subbytes_1_io_ret_1_3;
  wire       [7:0]    subbytes_1_io_ret_2_0;
  wire       [7:0]    subbytes_1_io_ret_2_1;
  wire       [7:0]    subbytes_1_io_ret_2_2;
  wire       [7:0]    subbytes_1_io_ret_2_3;
  wire       [7:0]    subbytes_1_io_ret_3_0;
  wire       [7:0]    subbytes_1_io_ret_3_1;
  wire       [7:0]    subbytes_1_io_ret_3_2;
  wire       [7:0]    subbytes_1_io_ret_3_3;
  wire       [7:0]    shiftrows_1_io_ret_0_0;
  wire       [7:0]    shiftrows_1_io_ret_0_1;
  wire       [7:0]    shiftrows_1_io_ret_0_2;
  wire       [7:0]    shiftrows_1_io_ret_0_3;
  wire       [7:0]    shiftrows_1_io_ret_1_0;
  wire       [7:0]    shiftrows_1_io_ret_1_1;
  wire       [7:0]    shiftrows_1_io_ret_1_2;
  wire       [7:0]    shiftrows_1_io_ret_1_3;
  wire       [7:0]    shiftrows_1_io_ret_2_0;
  wire       [7:0]    shiftrows_1_io_ret_2_1;
  wire       [7:0]    shiftrows_1_io_ret_2_2;
  wire       [7:0]    shiftrows_1_io_ret_2_3;
  wire       [7:0]    shiftrows_1_io_ret_3_0;
  wire       [7:0]    shiftrows_1_io_ret_3_1;
  wire       [7:0]    shiftrows_1_io_ret_3_2;
  wire       [7:0]    shiftrows_1_io_ret_3_3;
  wire       [7:0]    mixcolumns_1_io_ret_0_0;
  wire       [7:0]    mixcolumns_1_io_ret_0_1;
  wire       [7:0]    mixcolumns_1_io_ret_0_2;
  wire       [7:0]    mixcolumns_1_io_ret_0_3;
  wire       [7:0]    mixcolumns_1_io_ret_1_0;
  wire       [7:0]    mixcolumns_1_io_ret_1_1;
  wire       [7:0]    mixcolumns_1_io_ret_1_2;
  wire       [7:0]    mixcolumns_1_io_ret_1_3;
  wire       [7:0]    mixcolumns_1_io_ret_2_0;
  wire       [7:0]    mixcolumns_1_io_ret_2_1;
  wire       [7:0]    mixcolumns_1_io_ret_2_2;
  wire       [7:0]    mixcolumns_1_io_ret_2_3;
  wire       [7:0]    mixcolumns_1_io_ret_3_0;
  wire       [7:0]    mixcolumns_1_io_ret_3_1;
  wire       [7:0]    mixcolumns_1_io_ret_3_2;
  wire       [7:0]    mixcolumns_1_io_ret_3_3;
  wire       [7:0]    keyschedule_1_io_ret_0_0;
  wire       [7:0]    keyschedule_1_io_ret_0_1;
  wire       [7:0]    keyschedule_1_io_ret_0_2;
  wire       [7:0]    keyschedule_1_io_ret_0_3;
  wire       [7:0]    keyschedule_1_io_ret_1_0;
  wire       [7:0]    keyschedule_1_io_ret_1_1;
  wire       [7:0]    keyschedule_1_io_ret_1_2;
  wire       [7:0]    keyschedule_1_io_ret_1_3;
  wire       [7:0]    keyschedule_1_io_ret_2_0;
  wire       [7:0]    keyschedule_1_io_ret_2_1;
  wire       [7:0]    keyschedule_1_io_ret_2_2;
  wire       [7:0]    keyschedule_1_io_ret_2_3;
  wire       [7:0]    keyschedule_1_io_ret_3_0;
  wire       [7:0]    keyschedule_1_io_ret_3_1;
  wire       [7:0]    keyschedule_1_io_ret_3_2;
  wire       [7:0]    keyschedule_1_io_ret_3_3;
  wire       [7:0]    nextrc_1_io_ret;
  wire       [3:0]    _zz_counter_valueNext;
  wire       [0:0]    _zz_counter_valueNext_1;
  wire       [7:0]    state0_0_0;
  wire       [7:0]    state0_0_1;
  wire       [7:0]    state0_0_2;
  wire       [7:0]    state0_0_3;
  wire       [7:0]    state0_1_0;
  wire       [7:0]    state0_1_1;
  wire       [7:0]    state0_1_2;
  wire       [7:0]    state0_1_3;
  wire       [7:0]    state0_2_0;
  wire       [7:0]    state0_2_1;
  wire       [7:0]    state0_2_2;
  wire       [7:0]    state0_2_3;
  wire       [7:0]    state0_3_0;
  wire       [7:0]    state0_3_1;
  wire       [7:0]    state0_3_2;
  wire       [7:0]    state0_3_3;
  reg        [7:0]    rounds_0_0;
  reg        [7:0]    rounds_0_1;
  reg        [7:0]    rounds_0_2;
  reg        [7:0]    rounds_0_3;
  reg        [7:0]    rounds_1_0;
  reg        [7:0]    rounds_1_1;
  reg        [7:0]    rounds_1_2;
  reg        [7:0]    rounds_1_3;
  reg        [7:0]    rounds_2_0;
  reg        [7:0]    rounds_2_1;
  reg        [7:0]    rounds_2_2;
  reg        [7:0]    rounds_2_3;
  reg        [7:0]    rounds_3_0;
  reg        [7:0]    rounds_3_1;
  reg        [7:0]    rounds_3_2;
  reg        [7:0]    rounds_3_3;
  reg        [7:0]    keys_0_0;
  reg        [7:0]    keys_0_1;
  reg        [7:0]    keys_0_2;
  reg        [7:0]    keys_0_3;
  reg        [7:0]    keys_1_0;
  reg        [7:0]    keys_1_1;
  reg        [7:0]    keys_1_2;
  reg        [7:0]    keys_1_3;
  reg        [7:0]    keys_2_0;
  reg        [7:0]    keys_2_1;
  reg        [7:0]    keys_2_2;
  reg        [7:0]    keys_2_3;
  reg        [7:0]    keys_3_0;
  reg        [7:0]    keys_3_1;
  reg        [7:0]    keys_3_2;
  reg        [7:0]    keys_3_3;
  reg        [7:0]    rcs;
  reg                 counter_willIncrement;
  wire                counter_willClear;
  reg        [3:0]    counter_valueNext;
  reg        [3:0]    counter_value;
  wire                counter_willOverflowIfInc;
  wire                counter_willOverflow;
  reg                 fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg        [1:0]    fsm_stateReg;
  reg        [1:0]    fsm_stateNext;
  reg                 io_reset_regNext;
  wire                when_AES_Round_l50;
  reg        [127:0]  _zz_io_ret;
  wire                when_StateMachine_l235;
  `ifndef SYNTHESIS
  reg [111:0] fsm_stateReg_string;
  reg [111:0] fsm_stateNext_string;
  `endif


  assign _zz_counter_valueNext_1 = counter_willIncrement;
  assign _zz_counter_valueNext = {3'd0, _zz_counter_valueNext_1};
  AddRoundKey addroundkey_1 (
    .io_rk_0_0     (addroundkey_1_io_rk_0_0[7:0]   ), //i
    .io_rk_0_1     (addroundkey_1_io_rk_0_1[7:0]   ), //i
    .io_rk_0_2     (addroundkey_1_io_rk_0_2[7:0]   ), //i
    .io_rk_0_3     (addroundkey_1_io_rk_0_3[7:0]   ), //i
    .io_rk_1_0     (addroundkey_1_io_rk_1_0[7:0]   ), //i
    .io_rk_1_1     (addroundkey_1_io_rk_1_1[7:0]   ), //i
    .io_rk_1_2     (addroundkey_1_io_rk_1_2[7:0]   ), //i
    .io_rk_1_3     (addroundkey_1_io_rk_1_3[7:0]   ), //i
    .io_rk_2_0     (addroundkey_1_io_rk_2_0[7:0]   ), //i
    .io_rk_2_1     (addroundkey_1_io_rk_2_1[7:0]   ), //i
    .io_rk_2_2     (addroundkey_1_io_rk_2_2[7:0]   ), //i
    .io_rk_2_3     (addroundkey_1_io_rk_2_3[7:0]   ), //i
    .io_rk_3_0     (addroundkey_1_io_rk_3_0[7:0]   ), //i
    .io_rk_3_1     (addroundkey_1_io_rk_3_1[7:0]   ), //i
    .io_rk_3_2     (addroundkey_1_io_rk_3_2[7:0]   ), //i
    .io_rk_3_3     (addroundkey_1_io_rk_3_3[7:0]   ), //i
    .io_s_0_0      (addroundkey_1_io_s_0_0[7:0]    ), //i
    .io_s_0_1      (addroundkey_1_io_s_0_1[7:0]    ), //i
    .io_s_0_2      (addroundkey_1_io_s_0_2[7:0]    ), //i
    .io_s_0_3      (addroundkey_1_io_s_0_3[7:0]    ), //i
    .io_s_1_0      (addroundkey_1_io_s_1_0[7:0]    ), //i
    .io_s_1_1      (addroundkey_1_io_s_1_1[7:0]    ), //i
    .io_s_1_2      (addroundkey_1_io_s_1_2[7:0]    ), //i
    .io_s_1_3      (addroundkey_1_io_s_1_3[7:0]    ), //i
    .io_s_2_0      (addroundkey_1_io_s_2_0[7:0]    ), //i
    .io_s_2_1      (addroundkey_1_io_s_2_1[7:0]    ), //i
    .io_s_2_2      (addroundkey_1_io_s_2_2[7:0]    ), //i
    .io_s_2_3      (addroundkey_1_io_s_2_3[7:0]    ), //i
    .io_s_3_0      (addroundkey_1_io_s_3_0[7:0]    ), //i
    .io_s_3_1      (addroundkey_1_io_s_3_1[7:0]    ), //i
    .io_s_3_2      (addroundkey_1_io_s_3_2[7:0]    ), //i
    .io_s_3_3      (addroundkey_1_io_s_3_3[7:0]    ), //i
    .io_ret_0_0    (addroundkey_1_io_ret_0_0[7:0]  ), //o
    .io_ret_0_1    (addroundkey_1_io_ret_0_1[7:0]  ), //o
    .io_ret_0_2    (addroundkey_1_io_ret_0_2[7:0]  ), //o
    .io_ret_0_3    (addroundkey_1_io_ret_0_3[7:0]  ), //o
    .io_ret_1_0    (addroundkey_1_io_ret_1_0[7:0]  ), //o
    .io_ret_1_1    (addroundkey_1_io_ret_1_1[7:0]  ), //o
    .io_ret_1_2    (addroundkey_1_io_ret_1_2[7:0]  ), //o
    .io_ret_1_3    (addroundkey_1_io_ret_1_3[7:0]  ), //o
    .io_ret_2_0    (addroundkey_1_io_ret_2_0[7:0]  ), //o
    .io_ret_2_1    (addroundkey_1_io_ret_2_1[7:0]  ), //o
    .io_ret_2_2    (addroundkey_1_io_ret_2_2[7:0]  ), //o
    .io_ret_2_3    (addroundkey_1_io_ret_2_3[7:0]  ), //o
    .io_ret_3_0    (addroundkey_1_io_ret_3_0[7:0]  ), //o
    .io_ret_3_1    (addroundkey_1_io_ret_3_1[7:0]  ), //o
    .io_ret_3_2    (addroundkey_1_io_ret_3_2[7:0]  ), //o
    .io_ret_3_3    (addroundkey_1_io_ret_3_3[7:0]  )  //o
  );
  SubBytes subbytes_1 (
    .io_state_0_0    (rounds_0_0[7:0]             ), //i
    .io_state_0_1    (rounds_0_1[7:0]             ), //i
    .io_state_0_2    (rounds_0_2[7:0]             ), //i
    .io_state_0_3    (rounds_0_3[7:0]             ), //i
    .io_state_1_0    (rounds_1_0[7:0]             ), //i
    .io_state_1_1    (rounds_1_1[7:0]             ), //i
    .io_state_1_2    (rounds_1_2[7:0]             ), //i
    .io_state_1_3    (rounds_1_3[7:0]             ), //i
    .io_state_2_0    (rounds_2_0[7:0]             ), //i
    .io_state_2_1    (rounds_2_1[7:0]             ), //i
    .io_state_2_2    (rounds_2_2[7:0]             ), //i
    .io_state_2_3    (rounds_2_3[7:0]             ), //i
    .io_state_3_0    (rounds_3_0[7:0]             ), //i
    .io_state_3_1    (rounds_3_1[7:0]             ), //i
    .io_state_3_2    (rounds_3_2[7:0]             ), //i
    .io_state_3_3    (rounds_3_3[7:0]             ), //i
    .io_ret_0_0      (subbytes_1_io_ret_0_0[7:0]  ), //o
    .io_ret_0_1      (subbytes_1_io_ret_0_1[7:0]  ), //o
    .io_ret_0_2      (subbytes_1_io_ret_0_2[7:0]  ), //o
    .io_ret_0_3      (subbytes_1_io_ret_0_3[7:0]  ), //o
    .io_ret_1_0      (subbytes_1_io_ret_1_0[7:0]  ), //o
    .io_ret_1_1      (subbytes_1_io_ret_1_1[7:0]  ), //o
    .io_ret_1_2      (subbytes_1_io_ret_1_2[7:0]  ), //o
    .io_ret_1_3      (subbytes_1_io_ret_1_3[7:0]  ), //o
    .io_ret_2_0      (subbytes_1_io_ret_2_0[7:0]  ), //o
    .io_ret_2_1      (subbytes_1_io_ret_2_1[7:0]  ), //o
    .io_ret_2_2      (subbytes_1_io_ret_2_2[7:0]  ), //o
    .io_ret_2_3      (subbytes_1_io_ret_2_3[7:0]  ), //o
    .io_ret_3_0      (subbytes_1_io_ret_3_0[7:0]  ), //o
    .io_ret_3_1      (subbytes_1_io_ret_3_1[7:0]  ), //o
    .io_ret_3_2      (subbytes_1_io_ret_3_2[7:0]  ), //o
    .io_ret_3_3      (subbytes_1_io_ret_3_3[7:0]  )  //o
  );
  ShiftRows shiftrows_1 (
    .io_state_0_0    (subbytes_1_io_ret_0_0[7:0]   ), //i
    .io_state_0_1    (subbytes_1_io_ret_0_1[7:0]   ), //i
    .io_state_0_2    (subbytes_1_io_ret_0_2[7:0]   ), //i
    .io_state_0_3    (subbytes_1_io_ret_0_3[7:0]   ), //i
    .io_state_1_0    (subbytes_1_io_ret_1_0[7:0]   ), //i
    .io_state_1_1    (subbytes_1_io_ret_1_1[7:0]   ), //i
    .io_state_1_2    (subbytes_1_io_ret_1_2[7:0]   ), //i
    .io_state_1_3    (subbytes_1_io_ret_1_3[7:0]   ), //i
    .io_state_2_0    (subbytes_1_io_ret_2_0[7:0]   ), //i
    .io_state_2_1    (subbytes_1_io_ret_2_1[7:0]   ), //i
    .io_state_2_2    (subbytes_1_io_ret_2_2[7:0]   ), //i
    .io_state_2_3    (subbytes_1_io_ret_2_3[7:0]   ), //i
    .io_state_3_0    (subbytes_1_io_ret_3_0[7:0]   ), //i
    .io_state_3_1    (subbytes_1_io_ret_3_1[7:0]   ), //i
    .io_state_3_2    (subbytes_1_io_ret_3_2[7:0]   ), //i
    .io_state_3_3    (subbytes_1_io_ret_3_3[7:0]   ), //i
    .io_ret_0_0      (shiftrows_1_io_ret_0_0[7:0]  ), //o
    .io_ret_0_1      (shiftrows_1_io_ret_0_1[7:0]  ), //o
    .io_ret_0_2      (shiftrows_1_io_ret_0_2[7:0]  ), //o
    .io_ret_0_3      (shiftrows_1_io_ret_0_3[7:0]  ), //o
    .io_ret_1_0      (shiftrows_1_io_ret_1_0[7:0]  ), //o
    .io_ret_1_1      (shiftrows_1_io_ret_1_1[7:0]  ), //o
    .io_ret_1_2      (shiftrows_1_io_ret_1_2[7:0]  ), //o
    .io_ret_1_3      (shiftrows_1_io_ret_1_3[7:0]  ), //o
    .io_ret_2_0      (shiftrows_1_io_ret_2_0[7:0]  ), //o
    .io_ret_2_1      (shiftrows_1_io_ret_2_1[7:0]  ), //o
    .io_ret_2_2      (shiftrows_1_io_ret_2_2[7:0]  ), //o
    .io_ret_2_3      (shiftrows_1_io_ret_2_3[7:0]  ), //o
    .io_ret_3_0      (shiftrows_1_io_ret_3_0[7:0]  ), //o
    .io_ret_3_1      (shiftrows_1_io_ret_3_1[7:0]  ), //o
    .io_ret_3_2      (shiftrows_1_io_ret_3_2[7:0]  ), //o
    .io_ret_3_3      (shiftrows_1_io_ret_3_3[7:0]  )  //o
  );
  MixColumns mixcolumns_1 (
    .io_state_0_0    (shiftrows_1_io_ret_0_0[7:0]   ), //i
    .io_state_0_1    (shiftrows_1_io_ret_0_1[7:0]   ), //i
    .io_state_0_2    (shiftrows_1_io_ret_0_2[7:0]   ), //i
    .io_state_0_3    (shiftrows_1_io_ret_0_3[7:0]   ), //i
    .io_state_1_0    (shiftrows_1_io_ret_1_0[7:0]   ), //i
    .io_state_1_1    (shiftrows_1_io_ret_1_1[7:0]   ), //i
    .io_state_1_2    (shiftrows_1_io_ret_1_2[7:0]   ), //i
    .io_state_1_3    (shiftrows_1_io_ret_1_3[7:0]   ), //i
    .io_state_2_0    (shiftrows_1_io_ret_2_0[7:0]   ), //i
    .io_state_2_1    (shiftrows_1_io_ret_2_1[7:0]   ), //i
    .io_state_2_2    (shiftrows_1_io_ret_2_2[7:0]   ), //i
    .io_state_2_3    (shiftrows_1_io_ret_2_3[7:0]   ), //i
    .io_state_3_0    (shiftrows_1_io_ret_3_0[7:0]   ), //i
    .io_state_3_1    (shiftrows_1_io_ret_3_1[7:0]   ), //i
    .io_state_3_2    (shiftrows_1_io_ret_3_2[7:0]   ), //i
    .io_state_3_3    (shiftrows_1_io_ret_3_3[7:0]   ), //i
    .io_ret_0_0      (mixcolumns_1_io_ret_0_0[7:0]  ), //o
    .io_ret_0_1      (mixcolumns_1_io_ret_0_1[7:0]  ), //o
    .io_ret_0_2      (mixcolumns_1_io_ret_0_2[7:0]  ), //o
    .io_ret_0_3      (mixcolumns_1_io_ret_0_3[7:0]  ), //o
    .io_ret_1_0      (mixcolumns_1_io_ret_1_0[7:0]  ), //o
    .io_ret_1_1      (mixcolumns_1_io_ret_1_1[7:0]  ), //o
    .io_ret_1_2      (mixcolumns_1_io_ret_1_2[7:0]  ), //o
    .io_ret_1_3      (mixcolumns_1_io_ret_1_3[7:0]  ), //o
    .io_ret_2_0      (mixcolumns_1_io_ret_2_0[7:0]  ), //o
    .io_ret_2_1      (mixcolumns_1_io_ret_2_1[7:0]  ), //o
    .io_ret_2_2      (mixcolumns_1_io_ret_2_2[7:0]  ), //o
    .io_ret_2_3      (mixcolumns_1_io_ret_2_3[7:0]  ), //o
    .io_ret_3_0      (mixcolumns_1_io_ret_3_0[7:0]  ), //o
    .io_ret_3_1      (mixcolumns_1_io_ret_3_1[7:0]  ), //o
    .io_ret_3_2      (mixcolumns_1_io_ret_3_2[7:0]  ), //o
    .io_ret_3_3      (mixcolumns_1_io_ret_3_3[7:0]  )  //o
  );
  KeySchedule keyschedule_1 (
    .io_key_0_0    (keyschedule_1_io_key_0_0[7:0]  ), //i
    .io_key_0_1    (keyschedule_1_io_key_0_1[7:0]  ), //i
    .io_key_0_2    (keyschedule_1_io_key_0_2[7:0]  ), //i
    .io_key_0_3    (keyschedule_1_io_key_0_3[7:0]  ), //i
    .io_key_1_0    (keyschedule_1_io_key_1_0[7:0]  ), //i
    .io_key_1_1    (keyschedule_1_io_key_1_1[7:0]  ), //i
    .io_key_1_2    (keyschedule_1_io_key_1_2[7:0]  ), //i
    .io_key_1_3    (keyschedule_1_io_key_1_3[7:0]  ), //i
    .io_key_2_0    (keyschedule_1_io_key_2_0[7:0]  ), //i
    .io_key_2_1    (keyschedule_1_io_key_2_1[7:0]  ), //i
    .io_key_2_2    (keyschedule_1_io_key_2_2[7:0]  ), //i
    .io_key_2_3    (keyschedule_1_io_key_2_3[7:0]  ), //i
    .io_key_3_0    (keyschedule_1_io_key_3_0[7:0]  ), //i
    .io_key_3_1    (keyschedule_1_io_key_3_1[7:0]  ), //i
    .io_key_3_2    (keyschedule_1_io_key_3_2[7:0]  ), //i
    .io_key_3_3    (keyschedule_1_io_key_3_3[7:0]  ), //i
    .io_c          (rcs[7:0]                       ), //i
    .io_ret_0_0    (keyschedule_1_io_ret_0_0[7:0]  ), //o
    .io_ret_0_1    (keyschedule_1_io_ret_0_1[7:0]  ), //o
    .io_ret_0_2    (keyschedule_1_io_ret_0_2[7:0]  ), //o
    .io_ret_0_3    (keyschedule_1_io_ret_0_3[7:0]  ), //o
    .io_ret_1_0    (keyschedule_1_io_ret_1_0[7:0]  ), //o
    .io_ret_1_1    (keyschedule_1_io_ret_1_1[7:0]  ), //o
    .io_ret_1_2    (keyschedule_1_io_ret_1_2[7:0]  ), //o
    .io_ret_1_3    (keyschedule_1_io_ret_1_3[7:0]  ), //o
    .io_ret_2_0    (keyschedule_1_io_ret_2_0[7:0]  ), //o
    .io_ret_2_1    (keyschedule_1_io_ret_2_1[7:0]  ), //o
    .io_ret_2_2    (keyschedule_1_io_ret_2_2[7:0]  ), //o
    .io_ret_2_3    (keyschedule_1_io_ret_2_3[7:0]  ), //o
    .io_ret_3_0    (keyschedule_1_io_ret_3_0[7:0]  ), //o
    .io_ret_3_1    (keyschedule_1_io_ret_3_1[7:0]  ), //o
    .io_ret_3_2    (keyschedule_1_io_ret_3_2[7:0]  ), //o
    .io_ret_3_3    (keyschedule_1_io_ret_3_3[7:0]  )  //o
  );
  NextRC nextrc_1 (
    .io_rc     (rcs[7:0]              ), //i
    .io_ret    (nextrc_1_io_ret[7:0]  )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_BOOT : fsm_stateReg_string = "BOOT          ";
      fsm_enumDef_sReset : fsm_stateReg_string = "sReset        ";
      fsm_enumDef_sAESRound : fsm_stateReg_string = "sAESRound     ";
      fsm_enumDef_sAESFinalRound : fsm_stateReg_string = "sAESFinalRound";
      default : fsm_stateReg_string = "??????????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_BOOT : fsm_stateNext_string = "BOOT          ";
      fsm_enumDef_sReset : fsm_stateNext_string = "sReset        ";
      fsm_enumDef_sAESRound : fsm_stateNext_string = "sAESRound     ";
      fsm_enumDef_sAESFinalRound : fsm_stateNext_string = "sAESFinalRound";
      default : fsm_stateNext_string = "??????????????";
    endcase
  end
  `endif

  always @(*) begin
    counter_willIncrement = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
      end
      fsm_enumDef_sAESRound : begin
        counter_willIncrement = 1'b1;
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  assign counter_willClear = 1'b0;
  assign counter_willOverflowIfInc = (counter_value == 4'b1000);
  assign counter_willOverflow = (counter_willOverflowIfInc && counter_willIncrement);
  always @(*) begin
    if(counter_willOverflow) begin
      counter_valueNext = 4'b0000;
    end else begin
      counter_valueNext = (counter_value + _zz_counter_valueNext);
    end
    if(counter_willClear) begin
      counter_valueNext = 4'b0000;
    end
  end

  always @(*) begin
    io_ret = 128'h0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        io_ret = _zz_io_ret;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_done = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        io_done = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_0_0 = mixcolumns_1_io_ret_0_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_0_0 = io_pt[127 : 120];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_0_0 = shiftrows_1_io_ret_0_0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_0_1 = mixcolumns_1_io_ret_0_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_0_1 = io_pt[95 : 88];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_0_1 = shiftrows_1_io_ret_0_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_0_2 = mixcolumns_1_io_ret_0_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_0_2 = io_pt[63 : 56];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_0_2 = shiftrows_1_io_ret_0_2;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_0_3 = mixcolumns_1_io_ret_0_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_0_3 = io_pt[31 : 24];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_0_3 = shiftrows_1_io_ret_0_3;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_1_0 = mixcolumns_1_io_ret_1_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_1_0 = io_pt[119 : 112];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_1_0 = shiftrows_1_io_ret_1_0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_1_1 = mixcolumns_1_io_ret_1_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_1_1 = io_pt[87 : 80];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_1_1 = shiftrows_1_io_ret_1_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_1_2 = mixcolumns_1_io_ret_1_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_1_2 = io_pt[55 : 48];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_1_2 = shiftrows_1_io_ret_1_2;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_1_3 = mixcolumns_1_io_ret_1_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_1_3 = io_pt[23 : 16];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_1_3 = shiftrows_1_io_ret_1_3;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_2_0 = mixcolumns_1_io_ret_2_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_2_0 = io_pt[111 : 104];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_2_0 = shiftrows_1_io_ret_2_0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_2_1 = mixcolumns_1_io_ret_2_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_2_1 = io_pt[79 : 72];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_2_1 = shiftrows_1_io_ret_2_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_2_2 = mixcolumns_1_io_ret_2_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_2_2 = io_pt[47 : 40];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_2_2 = shiftrows_1_io_ret_2_2;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_2_3 = mixcolumns_1_io_ret_2_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_2_3 = io_pt[15 : 8];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_2_3 = shiftrows_1_io_ret_2_3;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_3_0 = mixcolumns_1_io_ret_3_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_3_0 = io_pt[103 : 96];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_3_0 = shiftrows_1_io_ret_3_0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_3_1 = mixcolumns_1_io_ret_3_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_3_1 = io_pt[71 : 64];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_3_1 = shiftrows_1_io_ret_3_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_3_2 = mixcolumns_1_io_ret_3_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_3_2 = io_pt[39 : 32];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_3_2 = shiftrows_1_io_ret_3_2;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_s_3_3 = mixcolumns_1_io_ret_3_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_s_3_3 = io_pt[7 : 0];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        addroundkey_1_io_s_3_3 = shiftrows_1_io_ret_3_3;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_0_0 = keys_0_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_0_0 = io_key[127 : 120];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_0_1 = keys_0_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_0_1 = io_key[95 : 88];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_0_2 = keys_0_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_0_2 = io_key[63 : 56];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_0_3 = keys_0_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_0_3 = io_key[31 : 24];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_1_0 = keys_1_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_1_0 = io_key[119 : 112];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_1_1 = keys_1_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_1_1 = io_key[87 : 80];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_1_2 = keys_1_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_1_2 = io_key[55 : 48];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_1_3 = keys_1_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_1_3 = io_key[23 : 16];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_2_0 = keys_2_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_2_0 = io_key[111 : 104];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_2_1 = keys_2_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_2_1 = io_key[79 : 72];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_2_2 = keys_2_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_2_2 = io_key[47 : 40];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_2_3 = keys_2_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_2_3 = io_key[15 : 8];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_3_0 = keys_3_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_3_0 = io_key[103 : 96];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_3_1 = keys_3_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_3_1 = io_key[71 : 64];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_3_2 = keys_3_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_3_2 = io_key[39 : 32];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    addroundkey_1_io_rk_3_3 = keys_3_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          addroundkey_1_io_rk_3_3 = io_key[7 : 0];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  assign state0_0_0 = addroundkey_1_io_ret_0_0;
  assign state0_0_1 = addroundkey_1_io_ret_0_1;
  assign state0_0_2 = addroundkey_1_io_ret_0_2;
  assign state0_0_3 = addroundkey_1_io_ret_0_3;
  assign state0_1_0 = addroundkey_1_io_ret_1_0;
  assign state0_1_1 = addroundkey_1_io_ret_1_1;
  assign state0_1_2 = addroundkey_1_io_ret_1_2;
  assign state0_1_3 = addroundkey_1_io_ret_1_3;
  assign state0_2_0 = addroundkey_1_io_ret_2_0;
  assign state0_2_1 = addroundkey_1_io_ret_2_1;
  assign state0_2_2 = addroundkey_1_io_ret_2_2;
  assign state0_2_3 = addroundkey_1_io_ret_2_3;
  assign state0_3_0 = addroundkey_1_io_ret_3_0;
  assign state0_3_1 = addroundkey_1_io_ret_3_1;
  assign state0_3_2 = addroundkey_1_io_ret_3_2;
  assign state0_3_3 = addroundkey_1_io_ret_3_3;
  always @(*) begin
    keyschedule_1_io_key_0_0 = keys_0_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_0_0 = io_key[127 : 120];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_0_1 = keys_0_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_0_1 = io_key[95 : 88];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_0_2 = keys_0_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_0_2 = io_key[63 : 56];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_0_3 = keys_0_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_0_3 = io_key[31 : 24];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_1_0 = keys_1_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_1_0 = io_key[119 : 112];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_1_1 = keys_1_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_1_1 = io_key[87 : 80];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_1_2 = keys_1_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_1_2 = io_key[55 : 48];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_1_3 = keys_1_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_1_3 = io_key[23 : 16];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_2_0 = keys_2_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_2_0 = io_key[111 : 104];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_2_1 = keys_2_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_2_1 = io_key[79 : 72];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_2_2 = keys_2_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_2_2 = io_key[47 : 40];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_2_3 = keys_2_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_2_3 = io_key[15 : 8];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_3_0 = keys_3_0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_3_0 = io_key[103 : 96];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_3_1 = keys_3_1;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_3_1 = io_key[71 : 64];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_3_2 = keys_3_2;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_3_2 = io_key[39 : 32];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    keyschedule_1_io_key_3_3 = keys_3_3;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          keyschedule_1_io_key_3_3 = io_key[7 : 0];
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fsm_wantExit = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
        fsm_wantExit = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          fsm_stateNext = fsm_enumDef_sAESRound;
        end
      end
      fsm_enumDef_sAESRound : begin
        if(counter_willOverflow) begin
          fsm_stateNext = fsm_enumDef_sAESFinalRound;
        end
      end
      fsm_enumDef_sAESFinalRound : begin
        fsm_stateNext = fsm_enumDef_BOOT;
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_enumDef_sReset;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_BOOT;
    end
  end

  assign when_AES_Round_l50 = ((! io_reset) && io_reset_regNext);
  always @(*) begin
    _zz_io_ret[127 : 120] = addroundkey_1_io_ret_0_0;
    _zz_io_ret[95 : 88] = addroundkey_1_io_ret_0_1;
    _zz_io_ret[63 : 56] = addroundkey_1_io_ret_0_2;
    _zz_io_ret[31 : 24] = addroundkey_1_io_ret_0_3;
    _zz_io_ret[119 : 112] = addroundkey_1_io_ret_1_0;
    _zz_io_ret[87 : 80] = addroundkey_1_io_ret_1_1;
    _zz_io_ret[55 : 48] = addroundkey_1_io_ret_1_2;
    _zz_io_ret[23 : 16] = addroundkey_1_io_ret_1_3;
    _zz_io_ret[111 : 104] = addroundkey_1_io_ret_2_0;
    _zz_io_ret[79 : 72] = addroundkey_1_io_ret_2_1;
    _zz_io_ret[47 : 40] = addroundkey_1_io_ret_2_2;
    _zz_io_ret[15 : 8] = addroundkey_1_io_ret_2_3;
    _zz_io_ret[103 : 96] = addroundkey_1_io_ret_3_0;
    _zz_io_ret[71 : 64] = addroundkey_1_io_ret_3_1;
    _zz_io_ret[39 : 32] = addroundkey_1_io_ret_3_2;
    _zz_io_ret[7 : 0] = addroundkey_1_io_ret_3_3;
  end

  assign when_StateMachine_l235 = ((! (fsm_stateReg == fsm_enumDef_sReset)) && (fsm_stateNext == fsm_enumDef_sReset));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      counter_value <= 4'b0000;
      fsm_stateReg <= fsm_enumDef_BOOT;
    end else begin
      counter_value <= counter_valueNext;
      fsm_stateReg <= fsm_stateNext;
    end
  end

  always @(posedge clk) begin
    rounds_0_0 <= addroundkey_1_io_ret_0_0;
    rounds_0_1 <= addroundkey_1_io_ret_0_1;
    rounds_0_2 <= addroundkey_1_io_ret_0_2;
    rounds_0_3 <= addroundkey_1_io_ret_0_3;
    rounds_1_0 <= addroundkey_1_io_ret_1_0;
    rounds_1_1 <= addroundkey_1_io_ret_1_1;
    rounds_1_2 <= addroundkey_1_io_ret_1_2;
    rounds_1_3 <= addroundkey_1_io_ret_1_3;
    rounds_2_0 <= addroundkey_1_io_ret_2_0;
    rounds_2_1 <= addroundkey_1_io_ret_2_1;
    rounds_2_2 <= addroundkey_1_io_ret_2_2;
    rounds_2_3 <= addroundkey_1_io_ret_2_3;
    rounds_3_0 <= addroundkey_1_io_ret_3_0;
    rounds_3_1 <= addroundkey_1_io_ret_3_1;
    rounds_3_2 <= addroundkey_1_io_ret_3_2;
    rounds_3_3 <= addroundkey_1_io_ret_3_3;
    keys_0_0 <= keyschedule_1_io_ret_0_0;
    keys_0_1 <= keyschedule_1_io_ret_0_1;
    keys_0_2 <= keyschedule_1_io_ret_0_2;
    keys_0_3 <= keyschedule_1_io_ret_0_3;
    keys_1_0 <= keyschedule_1_io_ret_1_0;
    keys_1_1 <= keyschedule_1_io_ret_1_1;
    keys_1_2 <= keyschedule_1_io_ret_1_2;
    keys_1_3 <= keyschedule_1_io_ret_1_3;
    keys_2_0 <= keyschedule_1_io_ret_2_0;
    keys_2_1 <= keyschedule_1_io_ret_2_1;
    keys_2_2 <= keyschedule_1_io_ret_2_2;
    keys_2_3 <= keyschedule_1_io_ret_2_3;
    keys_3_0 <= keyschedule_1_io_ret_3_0;
    keys_3_1 <= keyschedule_1_io_ret_3_1;
    keys_3_2 <= keyschedule_1_io_ret_3_2;
    keys_3_3 <= keyschedule_1_io_ret_3_3;
    rcs <= nextrc_1_io_ret;
    case(fsm_stateReg)
      fsm_enumDef_sReset : begin
        if(when_AES_Round_l50) begin
          rounds_0_0 <= state0_0_0;
          rounds_0_1 <= state0_0_1;
          rounds_0_2 <= state0_0_2;
          rounds_0_3 <= state0_0_3;
          rounds_1_0 <= state0_1_0;
          rounds_1_1 <= state0_1_1;
          rounds_1_2 <= state0_1_2;
          rounds_1_3 <= state0_1_3;
          rounds_2_0 <= state0_2_0;
          rounds_2_1 <= state0_2_1;
          rounds_2_2 <= state0_2_2;
          rounds_2_3 <= state0_2_3;
          rounds_3_0 <= state0_3_0;
          rounds_3_1 <= state0_3_1;
          rounds_3_2 <= state0_3_2;
          rounds_3_3 <= state0_3_3;
          rcs <= nextrc_1_io_ret;
        end
      end
      fsm_enumDef_sAESRound : begin
      end
      fsm_enumDef_sAESFinalRound : begin
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l235) begin
      rcs <= 8'h01;
    end
  end

  always @(posedge clk) begin
    io_reset_regNext <= io_reset;
  end


endmodule

module NextRC (
  input      [7:0]    io_rc,
  output reg [7:0]    io_ret
);

  wire       [7:0]    _zz_io_ret;
  wire                when_AES_Round_l196;

  assign _zz_io_ret = (io_rc <<< 1);
  assign when_AES_Round_l196 = (io_rc[7] == 1'b0);
  always @(*) begin
    if(when_AES_Round_l196) begin
      io_ret = (io_rc <<< 1);
    end else begin
      io_ret = (_zz_io_ret ^ 8'h1b);
    end
  end


endmodule

module KeySchedule (
  input      [7:0]    io_key_0_0,
  input      [7:0]    io_key_0_1,
  input      [7:0]    io_key_0_2,
  input      [7:0]    io_key_0_3,
  input      [7:0]    io_key_1_0,
  input      [7:0]    io_key_1_1,
  input      [7:0]    io_key_1_2,
  input      [7:0]    io_key_1_3,
  input      [7:0]    io_key_2_0,
  input      [7:0]    io_key_2_1,
  input      [7:0]    io_key_2_2,
  input      [7:0]    io_key_2_3,
  input      [7:0]    io_key_3_0,
  input      [7:0]    io_key_3_1,
  input      [7:0]    io_key_3_2,
  input      [7:0]    io_key_3_3,
  input      [7:0]    io_c,
  output     [7:0]    io_ret_0_0,
  output     [7:0]    io_ret_0_1,
  output     [7:0]    io_ret_0_2,
  output     [7:0]    io_ret_0_3,
  output     [7:0]    io_ret_1_0,
  output     [7:0]    io_ret_1_1,
  output     [7:0]    io_ret_1_2,
  output     [7:0]    io_ret_1_3,
  output     [7:0]    io_ret_2_0,
  output     [7:0]    io_ret_2_1,
  output     [7:0]    io_ret_2_2,
  output     [7:0]    io_ret_2_3,
  output     [7:0]    io_ret_3_0,
  output     [7:0]    io_ret_3_1,
  output     [7:0]    io_ret_3_2,
  output     [7:0]    io_ret_3_3
);

  wire       [7:0]    subword_1_io_ret_0;
  wire       [7:0]    subword_1_io_ret_1;
  wire       [7:0]    subword_1_io_ret_2;
  wire       [7:0]    subword_1_io_ret_3;
  wire       [7:0]    keyT_0_0;
  wire       [7:0]    keyT_0_1;
  wire       [7:0]    keyT_0_2;
  wire       [7:0]    keyT_0_3;
  wire       [7:0]    keyT_1_0;
  wire       [7:0]    keyT_1_1;
  wire       [7:0]    keyT_1_2;
  wire       [7:0]    keyT_1_3;
  wire       [7:0]    keyT_2_0;
  wire       [7:0]    keyT_2_1;
  wire       [7:0]    keyT_2_2;
  wire       [7:0]    keyT_2_3;
  wire       [7:0]    keyT_3_0;
  wire       [7:0]    keyT_3_1;
  wire       [7:0]    keyT_3_2;
  wire       [7:0]    keyT_3_3;
  wire       [7:0]    w0_0;
  wire       [7:0]    w0_1;
  wire       [7:0]    w0_2;
  wire       [7:0]    w0_3;
  wire       [7:0]    w1_0;
  wire       [7:0]    w1_1;
  wire       [7:0]    w1_2;
  wire       [7:0]    w1_3;
  wire       [7:0]    w2_0;
  wire       [7:0]    w2_1;
  wire       [7:0]    w2_2;
  wire       [7:0]    w2_3;
  wire       [7:0]    w3_0;
  wire       [7:0]    w3_1;
  wire       [7:0]    w3_2;
  wire       [7:0]    w3_3;

  SubWord subword_1 (
    .io_bs_0     (keyT_3_0[7:0]            ), //i
    .io_bs_1     (keyT_3_1[7:0]            ), //i
    .io_bs_2     (keyT_3_2[7:0]            ), //i
    .io_bs_3     (keyT_3_3[7:0]            ), //i
    .io_ret_0    (subword_1_io_ret_0[7:0]  ), //o
    .io_ret_1    (subword_1_io_ret_1[7:0]  ), //o
    .io_ret_2    (subword_1_io_ret_2[7:0]  ), //o
    .io_ret_3    (subword_1_io_ret_3[7:0]  )  //o
  );
  assign keyT_0_0 = io_key_0_0;
  assign keyT_0_1 = io_key_1_0;
  assign keyT_0_2 = io_key_2_0;
  assign keyT_0_3 = io_key_3_0;
  assign keyT_1_0 = io_key_0_1;
  assign keyT_1_1 = io_key_1_1;
  assign keyT_1_2 = io_key_2_1;
  assign keyT_1_3 = io_key_3_1;
  assign keyT_2_0 = io_key_0_2;
  assign keyT_2_1 = io_key_1_2;
  assign keyT_2_2 = io_key_2_2;
  assign keyT_2_3 = io_key_3_2;
  assign keyT_3_0 = io_key_0_3;
  assign keyT_3_1 = io_key_1_3;
  assign keyT_3_2 = io_key_2_3;
  assign keyT_3_3 = io_key_3_3;
  assign w0_0 = ((keyT_0_0 ^ subword_1_io_ret_1) ^ io_c);
  assign w0_1 = ((keyT_0_1 ^ subword_1_io_ret_2) ^ 8'h0);
  assign w0_2 = ((keyT_0_2 ^ subword_1_io_ret_3) ^ 8'h0);
  assign w0_3 = ((keyT_0_3 ^ subword_1_io_ret_0) ^ 8'h0);
  assign w1_0 = (keyT_1_0 ^ w0_0);
  assign w1_1 = (keyT_1_1 ^ w0_1);
  assign w1_2 = (keyT_1_2 ^ w0_2);
  assign w1_3 = (keyT_1_3 ^ w0_3);
  assign w2_0 = (keyT_2_0 ^ w1_0);
  assign w2_1 = (keyT_2_1 ^ w1_1);
  assign w2_2 = (keyT_2_2 ^ w1_2);
  assign w2_3 = (keyT_2_3 ^ w1_3);
  assign w3_0 = (keyT_3_0 ^ w2_0);
  assign w3_1 = (keyT_3_1 ^ w2_1);
  assign w3_2 = (keyT_3_2 ^ w2_2);
  assign w3_3 = (keyT_3_3 ^ w2_3);
  assign io_ret_0_0 = w0_0;
  assign io_ret_0_1 = w1_0;
  assign io_ret_0_2 = w2_0;
  assign io_ret_0_3 = w3_0;
  assign io_ret_1_0 = w0_1;
  assign io_ret_1_1 = w1_1;
  assign io_ret_1_2 = w2_1;
  assign io_ret_1_3 = w3_1;
  assign io_ret_2_0 = w0_2;
  assign io_ret_2_1 = w1_2;
  assign io_ret_2_2 = w2_2;
  assign io_ret_2_3 = w3_2;
  assign io_ret_3_0 = w0_3;
  assign io_ret_3_1 = w1_3;
  assign io_ret_3_2 = w2_3;
  assign io_ret_3_3 = w3_3;

endmodule

module MixColumns (
  input      [7:0]    io_state_0_0,
  input      [7:0]    io_state_0_1,
  input      [7:0]    io_state_0_2,
  input      [7:0]    io_state_0_3,
  input      [7:0]    io_state_1_0,
  input      [7:0]    io_state_1_1,
  input      [7:0]    io_state_1_2,
  input      [7:0]    io_state_1_3,
  input      [7:0]    io_state_2_0,
  input      [7:0]    io_state_2_1,
  input      [7:0]    io_state_2_2,
  input      [7:0]    io_state_2_3,
  input      [7:0]    io_state_3_0,
  input      [7:0]    io_state_3_1,
  input      [7:0]    io_state_3_2,
  input      [7:0]    io_state_3_3,
  output     [7:0]    io_ret_0_0,
  output     [7:0]    io_ret_0_1,
  output     [7:0]    io_ret_0_2,
  output     [7:0]    io_ret_0_3,
  output     [7:0]    io_ret_1_0,
  output     [7:0]    io_ret_1_1,
  output     [7:0]    io_ret_1_2,
  output     [7:0]    io_ret_1_3,
  output     [7:0]    io_ret_2_0,
  output     [7:0]    io_ret_2_1,
  output     [7:0]    io_ret_2_2,
  output     [7:0]    io_ret_2_3,
  output     [7:0]    io_ret_3_0,
  output     [7:0]    io_ret_3_1,
  output     [7:0]    io_ret_3_2,
  output     [7:0]    io_ret_3_3
);

  wire       [7:0]    mixColumn_4_io_ret_0;
  wire       [7:0]    mixColumn_4_io_ret_1;
  wire       [7:0]    mixColumn_4_io_ret_2;
  wire       [7:0]    mixColumn_4_io_ret_3;
  wire       [7:0]    mixColumn_5_io_ret_0;
  wire       [7:0]    mixColumn_5_io_ret_1;
  wire       [7:0]    mixColumn_5_io_ret_2;
  wire       [7:0]    mixColumn_5_io_ret_3;
  wire       [7:0]    mixColumn_6_io_ret_0;
  wire       [7:0]    mixColumn_6_io_ret_1;
  wire       [7:0]    mixColumn_6_io_ret_2;
  wire       [7:0]    mixColumn_6_io_ret_3;
  wire       [7:0]    mixColumn_7_io_ret_0;
  wire       [7:0]    mixColumn_7_io_ret_1;
  wire       [7:0]    mixColumn_7_io_ret_2;
  wire       [7:0]    mixColumn_7_io_ret_3;
  wire       [7:0]    ret_0_0;
  wire       [7:0]    ret_0_1;
  wire       [7:0]    ret_0_2;
  wire       [7:0]    ret_0_3;
  wire       [7:0]    ret_1_0;
  wire       [7:0]    ret_1_1;
  wire       [7:0]    ret_1_2;
  wire       [7:0]    ret_1_3;
  wire       [7:0]    ret_2_0;
  wire       [7:0]    ret_2_1;
  wire       [7:0]    ret_2_2;
  wire       [7:0]    ret_2_3;
  wire       [7:0]    ret_3_0;
  wire       [7:0]    ret_3_1;
  wire       [7:0]    ret_3_2;
  wire       [7:0]    ret_3_3;

  MixColumn mixColumn_4 (
    .io_c_0      (io_state_0_0[7:0]          ), //i
    .io_c_1      (io_state_1_0[7:0]          ), //i
    .io_c_2      (io_state_2_0[7:0]          ), //i
    .io_c_3      (io_state_3_0[7:0]          ), //i
    .io_ret_0    (mixColumn_4_io_ret_0[7:0]  ), //o
    .io_ret_1    (mixColumn_4_io_ret_1[7:0]  ), //o
    .io_ret_2    (mixColumn_4_io_ret_2[7:0]  ), //o
    .io_ret_3    (mixColumn_4_io_ret_3[7:0]  )  //o
  );
  MixColumn mixColumn_5 (
    .io_c_0      (io_state_0_1[7:0]          ), //i
    .io_c_1      (io_state_1_1[7:0]          ), //i
    .io_c_2      (io_state_2_1[7:0]          ), //i
    .io_c_3      (io_state_3_1[7:0]          ), //i
    .io_ret_0    (mixColumn_5_io_ret_0[7:0]  ), //o
    .io_ret_1    (mixColumn_5_io_ret_1[7:0]  ), //o
    .io_ret_2    (mixColumn_5_io_ret_2[7:0]  ), //o
    .io_ret_3    (mixColumn_5_io_ret_3[7:0]  )  //o
  );
  MixColumn mixColumn_6 (
    .io_c_0      (io_state_0_2[7:0]          ), //i
    .io_c_1      (io_state_1_2[7:0]          ), //i
    .io_c_2      (io_state_2_2[7:0]          ), //i
    .io_c_3      (io_state_3_2[7:0]          ), //i
    .io_ret_0    (mixColumn_6_io_ret_0[7:0]  ), //o
    .io_ret_1    (mixColumn_6_io_ret_1[7:0]  ), //o
    .io_ret_2    (mixColumn_6_io_ret_2[7:0]  ), //o
    .io_ret_3    (mixColumn_6_io_ret_3[7:0]  )  //o
  );
  MixColumn mixColumn_7 (
    .io_c_0      (io_state_0_3[7:0]          ), //i
    .io_c_1      (io_state_1_3[7:0]          ), //i
    .io_c_2      (io_state_2_3[7:0]          ), //i
    .io_c_3      (io_state_3_3[7:0]          ), //i
    .io_ret_0    (mixColumn_7_io_ret_0[7:0]  ), //o
    .io_ret_1    (mixColumn_7_io_ret_1[7:0]  ), //o
    .io_ret_2    (mixColumn_7_io_ret_2[7:0]  ), //o
    .io_ret_3    (mixColumn_7_io_ret_3[7:0]  )  //o
  );
  assign ret_0_0 = mixColumn_4_io_ret_0;
  assign ret_0_1 = mixColumn_4_io_ret_1;
  assign ret_0_2 = mixColumn_4_io_ret_2;
  assign ret_0_3 = mixColumn_4_io_ret_3;
  assign ret_1_0 = mixColumn_5_io_ret_0;
  assign ret_1_1 = mixColumn_5_io_ret_1;
  assign ret_1_2 = mixColumn_5_io_ret_2;
  assign ret_1_3 = mixColumn_5_io_ret_3;
  assign ret_2_0 = mixColumn_6_io_ret_0;
  assign ret_2_1 = mixColumn_6_io_ret_1;
  assign ret_2_2 = mixColumn_6_io_ret_2;
  assign ret_2_3 = mixColumn_6_io_ret_3;
  assign ret_3_0 = mixColumn_7_io_ret_0;
  assign ret_3_1 = mixColumn_7_io_ret_1;
  assign ret_3_2 = mixColumn_7_io_ret_2;
  assign ret_3_3 = mixColumn_7_io_ret_3;
  assign io_ret_0_0 = ret_0_0;
  assign io_ret_0_1 = ret_1_0;
  assign io_ret_0_2 = ret_2_0;
  assign io_ret_0_3 = ret_3_0;
  assign io_ret_1_0 = ret_0_1;
  assign io_ret_1_1 = ret_1_1;
  assign io_ret_1_2 = ret_2_1;
  assign io_ret_1_3 = ret_3_1;
  assign io_ret_2_0 = ret_0_2;
  assign io_ret_2_1 = ret_1_2;
  assign io_ret_2_2 = ret_2_2;
  assign io_ret_2_3 = ret_3_2;
  assign io_ret_3_0 = ret_0_3;
  assign io_ret_3_1 = ret_1_3;
  assign io_ret_3_2 = ret_2_3;
  assign io_ret_3_3 = ret_3_3;

endmodule

module ShiftRows (
  input      [7:0]    io_state_0_0,
  input      [7:0]    io_state_0_1,
  input      [7:0]    io_state_0_2,
  input      [7:0]    io_state_0_3,
  input      [7:0]    io_state_1_0,
  input      [7:0]    io_state_1_1,
  input      [7:0]    io_state_1_2,
  input      [7:0]    io_state_1_3,
  input      [7:0]    io_state_2_0,
  input      [7:0]    io_state_2_1,
  input      [7:0]    io_state_2_2,
  input      [7:0]    io_state_2_3,
  input      [7:0]    io_state_3_0,
  input      [7:0]    io_state_3_1,
  input      [7:0]    io_state_3_2,
  input      [7:0]    io_state_3_3,
  output     [7:0]    io_ret_0_0,
  output     [7:0]    io_ret_0_1,
  output     [7:0]    io_ret_0_2,
  output     [7:0]    io_ret_0_3,
  output     [7:0]    io_ret_1_0,
  output     [7:0]    io_ret_1_1,
  output     [7:0]    io_ret_1_2,
  output     [7:0]    io_ret_1_3,
  output     [7:0]    io_ret_2_0,
  output     [7:0]    io_ret_2_1,
  output     [7:0]    io_ret_2_2,
  output     [7:0]    io_ret_2_3,
  output     [7:0]    io_ret_3_0,
  output     [7:0]    io_ret_3_1,
  output     [7:0]    io_ret_3_2,
  output     [7:0]    io_ret_3_3
);


  assign io_ret_0_0 = io_state_0_0;
  assign io_ret_0_1 = io_state_0_1;
  assign io_ret_0_2 = io_state_0_2;
  assign io_ret_0_3 = io_state_0_3;
  assign io_ret_1_0 = io_state_1_1;
  assign io_ret_1_1 = io_state_1_2;
  assign io_ret_1_2 = io_state_1_3;
  assign io_ret_1_3 = io_state_1_0;
  assign io_ret_2_0 = io_state_2_2;
  assign io_ret_2_1 = io_state_2_3;
  assign io_ret_2_2 = io_state_2_0;
  assign io_ret_2_3 = io_state_2_1;
  assign io_ret_3_0 = io_state_3_3;
  assign io_ret_3_1 = io_state_3_0;
  assign io_ret_3_2 = io_state_3_1;
  assign io_ret_3_3 = io_state_3_2;

endmodule

module SubBytes (
  input      [7:0]    io_state_0_0,
  input      [7:0]    io_state_0_1,
  input      [7:0]    io_state_0_2,
  input      [7:0]    io_state_0_3,
  input      [7:0]    io_state_1_0,
  input      [7:0]    io_state_1_1,
  input      [7:0]    io_state_1_2,
  input      [7:0]    io_state_1_3,
  input      [7:0]    io_state_2_0,
  input      [7:0]    io_state_2_1,
  input      [7:0]    io_state_2_2,
  input      [7:0]    io_state_2_3,
  input      [7:0]    io_state_3_0,
  input      [7:0]    io_state_3_1,
  input      [7:0]    io_state_3_2,
  input      [7:0]    io_state_3_3,
  output     [7:0]    io_ret_0_0,
  output     [7:0]    io_ret_0_1,
  output     [7:0]    io_ret_0_2,
  output     [7:0]    io_ret_0_3,
  output     [7:0]    io_ret_1_0,
  output     [7:0]    io_ret_1_1,
  output     [7:0]    io_ret_1_2,
  output     [7:0]    io_ret_1_3,
  output     [7:0]    io_ret_2_0,
  output     [7:0]    io_ret_2_1,
  output     [7:0]    io_ret_2_2,
  output     [7:0]    io_ret_2_3,
  output     [7:0]    io_ret_3_0,
  output     [7:0]    io_ret_3_1,
  output     [7:0]    io_ret_3_2,
  output     [7:0]    io_ret_3_3
);

  wire       [7:0]    subByte_20_io_ret;
  wire       [7:0]    subByte_21_io_ret;
  wire       [7:0]    subByte_22_io_ret;
  wire       [7:0]    subByte_23_io_ret;
  wire       [7:0]    subByte_24_io_ret;
  wire       [7:0]    subByte_25_io_ret;
  wire       [7:0]    subByte_26_io_ret;
  wire       [7:0]    subByte_27_io_ret;
  wire       [7:0]    subByte_28_io_ret;
  wire       [7:0]    subByte_29_io_ret;
  wire       [7:0]    subByte_30_io_ret;
  wire       [7:0]    subByte_31_io_ret;
  wire       [7:0]    subByte_32_io_ret;
  wire       [7:0]    subByte_33_io_ret;
  wire       [7:0]    subByte_34_io_ret;
  wire       [7:0]    subByte_35_io_ret;

  SubByte subByte_20 (
    .io_b      (io_state_0_0[7:0]       ), //i
    .io_ret    (subByte_20_io_ret[7:0]  )  //o
  );
  SubByte subByte_21 (
    .io_b      (io_state_0_1[7:0]       ), //i
    .io_ret    (subByte_21_io_ret[7:0]  )  //o
  );
  SubByte subByte_22 (
    .io_b      (io_state_0_2[7:0]       ), //i
    .io_ret    (subByte_22_io_ret[7:0]  )  //o
  );
  SubByte subByte_23 (
    .io_b      (io_state_0_3[7:0]       ), //i
    .io_ret    (subByte_23_io_ret[7:0]  )  //o
  );
  SubByte subByte_24 (
    .io_b      (io_state_1_0[7:0]       ), //i
    .io_ret    (subByte_24_io_ret[7:0]  )  //o
  );
  SubByte subByte_25 (
    .io_b      (io_state_1_1[7:0]       ), //i
    .io_ret    (subByte_25_io_ret[7:0]  )  //o
  );
  SubByte subByte_26 (
    .io_b      (io_state_1_2[7:0]       ), //i
    .io_ret    (subByte_26_io_ret[7:0]  )  //o
  );
  SubByte subByte_27 (
    .io_b      (io_state_1_3[7:0]       ), //i
    .io_ret    (subByte_27_io_ret[7:0]  )  //o
  );
  SubByte subByte_28 (
    .io_b      (io_state_2_0[7:0]       ), //i
    .io_ret    (subByte_28_io_ret[7:0]  )  //o
  );
  SubByte subByte_29 (
    .io_b      (io_state_2_1[7:0]       ), //i
    .io_ret    (subByte_29_io_ret[7:0]  )  //o
  );
  SubByte subByte_30 (
    .io_b      (io_state_2_2[7:0]       ), //i
    .io_ret    (subByte_30_io_ret[7:0]  )  //o
  );
  SubByte subByte_31 (
    .io_b      (io_state_2_3[7:0]       ), //i
    .io_ret    (subByte_31_io_ret[7:0]  )  //o
  );
  SubByte subByte_32 (
    .io_b      (io_state_3_0[7:0]       ), //i
    .io_ret    (subByte_32_io_ret[7:0]  )  //o
  );
  SubByte subByte_33 (
    .io_b      (io_state_3_1[7:0]       ), //i
    .io_ret    (subByte_33_io_ret[7:0]  )  //o
  );
  SubByte subByte_34 (
    .io_b      (io_state_3_2[7:0]       ), //i
    .io_ret    (subByte_34_io_ret[7:0]  )  //o
  );
  SubByte subByte_35 (
    .io_b      (io_state_3_3[7:0]       ), //i
    .io_ret    (subByte_35_io_ret[7:0]  )  //o
  );
  assign io_ret_0_0 = subByte_20_io_ret;
  assign io_ret_0_1 = subByte_21_io_ret;
  assign io_ret_0_2 = subByte_22_io_ret;
  assign io_ret_0_3 = subByte_23_io_ret;
  assign io_ret_1_0 = subByte_24_io_ret;
  assign io_ret_1_1 = subByte_25_io_ret;
  assign io_ret_1_2 = subByte_26_io_ret;
  assign io_ret_1_3 = subByte_27_io_ret;
  assign io_ret_2_0 = subByte_28_io_ret;
  assign io_ret_2_1 = subByte_29_io_ret;
  assign io_ret_2_2 = subByte_30_io_ret;
  assign io_ret_2_3 = subByte_31_io_ret;
  assign io_ret_3_0 = subByte_32_io_ret;
  assign io_ret_3_1 = subByte_33_io_ret;
  assign io_ret_3_2 = subByte_34_io_ret;
  assign io_ret_3_3 = subByte_35_io_ret;

endmodule

module AddRoundKey (
  input      [7:0]    io_rk_0_0,
  input      [7:0]    io_rk_0_1,
  input      [7:0]    io_rk_0_2,
  input      [7:0]    io_rk_0_3,
  input      [7:0]    io_rk_1_0,
  input      [7:0]    io_rk_1_1,
  input      [7:0]    io_rk_1_2,
  input      [7:0]    io_rk_1_3,
  input      [7:0]    io_rk_2_0,
  input      [7:0]    io_rk_2_1,
  input      [7:0]    io_rk_2_2,
  input      [7:0]    io_rk_2_3,
  input      [7:0]    io_rk_3_0,
  input      [7:0]    io_rk_3_1,
  input      [7:0]    io_rk_3_2,
  input      [7:0]    io_rk_3_3,
  input      [7:0]    io_s_0_0,
  input      [7:0]    io_s_0_1,
  input      [7:0]    io_s_0_2,
  input      [7:0]    io_s_0_3,
  input      [7:0]    io_s_1_0,
  input      [7:0]    io_s_1_1,
  input      [7:0]    io_s_1_2,
  input      [7:0]    io_s_1_3,
  input      [7:0]    io_s_2_0,
  input      [7:0]    io_s_2_1,
  input      [7:0]    io_s_2_2,
  input      [7:0]    io_s_2_3,
  input      [7:0]    io_s_3_0,
  input      [7:0]    io_s_3_1,
  input      [7:0]    io_s_3_2,
  input      [7:0]    io_s_3_3,
  output     [7:0]    io_ret_0_0,
  output     [7:0]    io_ret_0_1,
  output     [7:0]    io_ret_0_2,
  output     [7:0]    io_ret_0_3,
  output     [7:0]    io_ret_1_0,
  output     [7:0]    io_ret_1_1,
  output     [7:0]    io_ret_1_2,
  output     [7:0]    io_ret_1_3,
  output     [7:0]    io_ret_2_0,
  output     [7:0]    io_ret_2_1,
  output     [7:0]    io_ret_2_2,
  output     [7:0]    io_ret_2_3,
  output     [7:0]    io_ret_3_0,
  output     [7:0]    io_ret_3_1,
  output     [7:0]    io_ret_3_2,
  output     [7:0]    io_ret_3_3
);


  assign io_ret_0_0 = (io_rk_0_0 ^ io_s_0_0);
  assign io_ret_0_1 = (io_rk_0_1 ^ io_s_0_1);
  assign io_ret_0_2 = (io_rk_0_2 ^ io_s_0_2);
  assign io_ret_0_3 = (io_rk_0_3 ^ io_s_0_3);
  assign io_ret_1_0 = (io_rk_1_0 ^ io_s_1_0);
  assign io_ret_1_1 = (io_rk_1_1 ^ io_s_1_1);
  assign io_ret_1_2 = (io_rk_1_2 ^ io_s_1_2);
  assign io_ret_1_3 = (io_rk_1_3 ^ io_s_1_3);
  assign io_ret_2_0 = (io_rk_2_0 ^ io_s_2_0);
  assign io_ret_2_1 = (io_rk_2_1 ^ io_s_2_1);
  assign io_ret_2_2 = (io_rk_2_2 ^ io_s_2_2);
  assign io_ret_2_3 = (io_rk_2_3 ^ io_s_2_3);
  assign io_ret_3_0 = (io_rk_3_0 ^ io_s_3_0);
  assign io_ret_3_1 = (io_rk_3_1 ^ io_s_3_1);
  assign io_ret_3_2 = (io_rk_3_2 ^ io_s_3_2);
  assign io_ret_3_3 = (io_rk_3_3 ^ io_s_3_3);

endmodule

module SubWord (
  input      [7:0]    io_bs_0,
  input      [7:0]    io_bs_1,
  input      [7:0]    io_bs_2,
  input      [7:0]    io_bs_3,
  output     [7:0]    io_ret_0,
  output     [7:0]    io_ret_1,
  output     [7:0]    io_ret_2,
  output     [7:0]    io_ret_3
);

  wire       [7:0]    subByte_20_io_ret;
  wire       [7:0]    subByte_21_io_ret;
  wire       [7:0]    subByte_22_io_ret;
  wire       [7:0]    subByte_23_io_ret;

  SubByte subByte_20 (
    .io_b      (io_bs_0[7:0]            ), //i
    .io_ret    (subByte_20_io_ret[7:0]  )  //o
  );
  SubByte subByte_21 (
    .io_b      (io_bs_1[7:0]            ), //i
    .io_ret    (subByte_21_io_ret[7:0]  )  //o
  );
  SubByte subByte_22 (
    .io_b      (io_bs_2[7:0]            ), //i
    .io_ret    (subByte_22_io_ret[7:0]  )  //o
  );
  SubByte subByte_23 (
    .io_b      (io_bs_3[7:0]            ), //i
    .io_ret    (subByte_23_io_ret[7:0]  )  //o
  );
  assign io_ret_0 = subByte_20_io_ret;
  assign io_ret_1 = subByte_21_io_ret;
  assign io_ret_2 = subByte_22_io_ret;
  assign io_ret_3 = subByte_23_io_ret;

endmodule

//MixColumn replaced by MixColumn

//MixColumn replaced by MixColumn

//MixColumn replaced by MixColumn

module MixColumn (
  input      [7:0]    io_c_0,
  input      [7:0]    io_c_1,
  input      [7:0]    io_c_2,
  input      [7:0]    io_c_3,
  output     [7:0]    io_ret_0,
  output     [7:0]    io_ret_1,
  output     [7:0]    io_ret_2,
  output     [7:0]    io_ret_3
);

  wire       [7:0]    _zz__zz_io_ret_0;
  wire       [7:0]    _zz__zz_io_ret_0_1;
  wire       [7:0]    _zz__zz_io_ret_1;
  wire       [7:0]    _zz__zz_io_ret_1_1;
  wire       [7:0]    _zz__zz_io_ret_2;
  wire       [7:0]    _zz__zz_io_ret_2_1;
  wire       [7:0]    _zz__zz_io_ret_3;
  wire       [7:0]    _zz__zz_io_ret_3_1;
  reg        [7:0]    _zz_io_ret_0;
  wire                when_AES_Round_l157;
  reg        [7:0]    _zz_io_ret_0_1;
  wire                when_AES_Round_l157_1;
  reg        [7:0]    _zz_io_ret_1;
  wire                when_AES_Round_l157_2;
  reg        [7:0]    _zz_io_ret_1_1;
  wire                when_AES_Round_l157_3;
  reg        [7:0]    _zz_io_ret_2;
  wire                when_AES_Round_l157_4;
  reg        [7:0]    _zz_io_ret_2_1;
  wire                when_AES_Round_l157_5;
  reg        [7:0]    _zz_io_ret_3;
  wire                when_AES_Round_l157_6;
  reg        [7:0]    _zz_io_ret_3_1;
  wire                when_AES_Round_l157_7;

  assign _zz__zz_io_ret_0 = (io_c_0 <<< 1);
  assign _zz__zz_io_ret_0_1 = (io_c_1 <<< 1);
  assign _zz__zz_io_ret_1 = (io_c_1 <<< 1);
  assign _zz__zz_io_ret_1_1 = (io_c_2 <<< 1);
  assign _zz__zz_io_ret_2 = (io_c_2 <<< 1);
  assign _zz__zz_io_ret_2_1 = (io_c_3 <<< 1);
  assign _zz__zz_io_ret_3 = (io_c_0 <<< 1);
  assign _zz__zz_io_ret_3_1 = (io_c_3 <<< 1);
  assign when_AES_Round_l157 = (io_c_0[7] == 1'b0);
  always @(*) begin
    if(when_AES_Round_l157) begin
      _zz_io_ret_0 = (io_c_0 <<< 1);
    end else begin
      _zz_io_ret_0 = (_zz__zz_io_ret_0 ^ 8'h1b);
    end
  end

  assign when_AES_Round_l157_1 = (io_c_1[7] == 1'b0);
  always @(*) begin
    if(when_AES_Round_l157_1) begin
      _zz_io_ret_0_1 = (io_c_1 <<< 1);
    end else begin
      _zz_io_ret_0_1 = (_zz__zz_io_ret_0_1 ^ 8'h1b);
    end
  end

  assign io_ret_0 = (((_zz_io_ret_0 ^ (_zz_io_ret_0_1 ^ io_c_1)) ^ io_c_2) ^ io_c_3);
  assign when_AES_Round_l157_2 = (io_c_1[7] == 1'b0);
  always @(*) begin
    if(when_AES_Round_l157_2) begin
      _zz_io_ret_1 = (io_c_1 <<< 1);
    end else begin
      _zz_io_ret_1 = (_zz__zz_io_ret_1 ^ 8'h1b);
    end
  end

  assign when_AES_Round_l157_3 = (io_c_2[7] == 1'b0);
  always @(*) begin
    if(when_AES_Round_l157_3) begin
      _zz_io_ret_1_1 = (io_c_2 <<< 1);
    end else begin
      _zz_io_ret_1_1 = (_zz__zz_io_ret_1_1 ^ 8'h1b);
    end
  end

  assign io_ret_1 = (((io_c_0 ^ _zz_io_ret_1) ^ (_zz_io_ret_1_1 ^ io_c_2)) ^ io_c_3);
  assign when_AES_Round_l157_4 = (io_c_2[7] == 1'b0);
  always @(*) begin
    if(when_AES_Round_l157_4) begin
      _zz_io_ret_2 = (io_c_2 <<< 1);
    end else begin
      _zz_io_ret_2 = (_zz__zz_io_ret_2 ^ 8'h1b);
    end
  end

  assign when_AES_Round_l157_5 = (io_c_3[7] == 1'b0);
  always @(*) begin
    if(when_AES_Round_l157_5) begin
      _zz_io_ret_2_1 = (io_c_3 <<< 1);
    end else begin
      _zz_io_ret_2_1 = (_zz__zz_io_ret_2_1 ^ 8'h1b);
    end
  end

  assign io_ret_2 = (((io_c_0 ^ io_c_1) ^ _zz_io_ret_2) ^ (_zz_io_ret_2_1 ^ io_c_3));
  assign when_AES_Round_l157_6 = (io_c_0[7] == 1'b0);
  always @(*) begin
    if(when_AES_Round_l157_6) begin
      _zz_io_ret_3 = (io_c_0 <<< 1);
    end else begin
      _zz_io_ret_3 = (_zz__zz_io_ret_3 ^ 8'h1b);
    end
  end

  assign when_AES_Round_l157_7 = (io_c_3[7] == 1'b0);
  always @(*) begin
    if(when_AES_Round_l157_7) begin
      _zz_io_ret_3_1 = (io_c_3 <<< 1);
    end else begin
      _zz_io_ret_3_1 = (_zz__zz_io_ret_3_1 ^ 8'h1b);
    end
  end

  assign io_ret_3 = ((((_zz_io_ret_3 ^ io_c_0) ^ io_c_1) ^ io_c_2) ^ _zz_io_ret_3_1);

endmodule

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

//SubByte replaced by SubByte

module SubByte (
  input      [7:0]    io_b,
  output     [7:0]    io_ret
);

  reg        [7:0]    _zz_io_ret;

  always @(*) begin
    case(io_b)
      8'h0 : begin
        _zz_io_ret = 8'h63;
      end
      8'h01 : begin
        _zz_io_ret = 8'h7c;
      end
      8'h02 : begin
        _zz_io_ret = 8'h77;
      end
      8'h03 : begin
        _zz_io_ret = 8'h7b;
      end
      8'h04 : begin
        _zz_io_ret = 8'hf2;
      end
      8'h05 : begin
        _zz_io_ret = 8'h6b;
      end
      8'h06 : begin
        _zz_io_ret = 8'h6f;
      end
      8'h07 : begin
        _zz_io_ret = 8'hc5;
      end
      8'h08 : begin
        _zz_io_ret = 8'h30;
      end
      8'h09 : begin
        _zz_io_ret = 8'h01;
      end
      8'h0a : begin
        _zz_io_ret = 8'h67;
      end
      8'h0b : begin
        _zz_io_ret = 8'h2b;
      end
      8'h0c : begin
        _zz_io_ret = 8'hfe;
      end
      8'h0d : begin
        _zz_io_ret = 8'hd7;
      end
      8'h0e : begin
        _zz_io_ret = 8'hab;
      end
      8'h0f : begin
        _zz_io_ret = 8'h76;
      end
      8'h10 : begin
        _zz_io_ret = 8'hca;
      end
      8'h11 : begin
        _zz_io_ret = 8'h82;
      end
      8'h12 : begin
        _zz_io_ret = 8'hc9;
      end
      8'h13 : begin
        _zz_io_ret = 8'h7d;
      end
      8'h14 : begin
        _zz_io_ret = 8'hfa;
      end
      8'h15 : begin
        _zz_io_ret = 8'h59;
      end
      8'h16 : begin
        _zz_io_ret = 8'h47;
      end
      8'h17 : begin
        _zz_io_ret = 8'hf0;
      end
      8'h18 : begin
        _zz_io_ret = 8'had;
      end
      8'h19 : begin
        _zz_io_ret = 8'hd4;
      end
      8'h1a : begin
        _zz_io_ret = 8'ha2;
      end
      8'h1b : begin
        _zz_io_ret = 8'haf;
      end
      8'h1c : begin
        _zz_io_ret = 8'h9c;
      end
      8'h1d : begin
        _zz_io_ret = 8'ha4;
      end
      8'h1e : begin
        _zz_io_ret = 8'h72;
      end
      8'h1f : begin
        _zz_io_ret = 8'hc0;
      end
      8'h20 : begin
        _zz_io_ret = 8'hb7;
      end
      8'h21 : begin
        _zz_io_ret = 8'hfd;
      end
      8'h22 : begin
        _zz_io_ret = 8'h93;
      end
      8'h23 : begin
        _zz_io_ret = 8'h26;
      end
      8'h24 : begin
        _zz_io_ret = 8'h36;
      end
      8'h25 : begin
        _zz_io_ret = 8'h3f;
      end
      8'h26 : begin
        _zz_io_ret = 8'hf7;
      end
      8'h27 : begin
        _zz_io_ret = 8'hcc;
      end
      8'h28 : begin
        _zz_io_ret = 8'h34;
      end
      8'h29 : begin
        _zz_io_ret = 8'ha5;
      end
      8'h2a : begin
        _zz_io_ret = 8'he5;
      end
      8'h2b : begin
        _zz_io_ret = 8'hf1;
      end
      8'h2c : begin
        _zz_io_ret = 8'h71;
      end
      8'h2d : begin
        _zz_io_ret = 8'hd8;
      end
      8'h2e : begin
        _zz_io_ret = 8'h31;
      end
      8'h2f : begin
        _zz_io_ret = 8'h15;
      end
      8'h30 : begin
        _zz_io_ret = 8'h04;
      end
      8'h31 : begin
        _zz_io_ret = 8'hc7;
      end
      8'h32 : begin
        _zz_io_ret = 8'h23;
      end
      8'h33 : begin
        _zz_io_ret = 8'hc3;
      end
      8'h34 : begin
        _zz_io_ret = 8'h18;
      end
      8'h35 : begin
        _zz_io_ret = 8'h96;
      end
      8'h36 : begin
        _zz_io_ret = 8'h05;
      end
      8'h37 : begin
        _zz_io_ret = 8'h9a;
      end
      8'h38 : begin
        _zz_io_ret = 8'h07;
      end
      8'h39 : begin
        _zz_io_ret = 8'h12;
      end
      8'h3a : begin
        _zz_io_ret = 8'h80;
      end
      8'h3b : begin
        _zz_io_ret = 8'he2;
      end
      8'h3c : begin
        _zz_io_ret = 8'heb;
      end
      8'h3d : begin
        _zz_io_ret = 8'h27;
      end
      8'h3e : begin
        _zz_io_ret = 8'hb2;
      end
      8'h3f : begin
        _zz_io_ret = 8'h75;
      end
      8'h40 : begin
        _zz_io_ret = 8'h09;
      end
      8'h41 : begin
        _zz_io_ret = 8'h83;
      end
      8'h42 : begin
        _zz_io_ret = 8'h2c;
      end
      8'h43 : begin
        _zz_io_ret = 8'h1a;
      end
      8'h44 : begin
        _zz_io_ret = 8'h1b;
      end
      8'h45 : begin
        _zz_io_ret = 8'h6e;
      end
      8'h46 : begin
        _zz_io_ret = 8'h5a;
      end
      8'h47 : begin
        _zz_io_ret = 8'ha0;
      end
      8'h48 : begin
        _zz_io_ret = 8'h52;
      end
      8'h49 : begin
        _zz_io_ret = 8'h3b;
      end
      8'h4a : begin
        _zz_io_ret = 8'hd6;
      end
      8'h4b : begin
        _zz_io_ret = 8'hb3;
      end
      8'h4c : begin
        _zz_io_ret = 8'h29;
      end
      8'h4d : begin
        _zz_io_ret = 8'he3;
      end
      8'h4e : begin
        _zz_io_ret = 8'h2f;
      end
      8'h4f : begin
        _zz_io_ret = 8'h84;
      end
      8'h50 : begin
        _zz_io_ret = 8'h53;
      end
      8'h51 : begin
        _zz_io_ret = 8'hd1;
      end
      8'h52 : begin
        _zz_io_ret = 8'h0;
      end
      8'h53 : begin
        _zz_io_ret = 8'hed;
      end
      8'h54 : begin
        _zz_io_ret = 8'h20;
      end
      8'h55 : begin
        _zz_io_ret = 8'hfc;
      end
      8'h56 : begin
        _zz_io_ret = 8'hb1;
      end
      8'h57 : begin
        _zz_io_ret = 8'h5b;
      end
      8'h58 : begin
        _zz_io_ret = 8'h6a;
      end
      8'h59 : begin
        _zz_io_ret = 8'hcb;
      end
      8'h5a : begin
        _zz_io_ret = 8'hbe;
      end
      8'h5b : begin
        _zz_io_ret = 8'h39;
      end
      8'h5c : begin
        _zz_io_ret = 8'h4a;
      end
      8'h5d : begin
        _zz_io_ret = 8'h4c;
      end
      8'h5e : begin
        _zz_io_ret = 8'h58;
      end
      8'h5f : begin
        _zz_io_ret = 8'hcf;
      end
      8'h60 : begin
        _zz_io_ret = 8'hd0;
      end
      8'h61 : begin
        _zz_io_ret = 8'hef;
      end
      8'h62 : begin
        _zz_io_ret = 8'haa;
      end
      8'h63 : begin
        _zz_io_ret = 8'hfb;
      end
      8'h64 : begin
        _zz_io_ret = 8'h43;
      end
      8'h65 : begin
        _zz_io_ret = 8'h4d;
      end
      8'h66 : begin
        _zz_io_ret = 8'h33;
      end
      8'h67 : begin
        _zz_io_ret = 8'h85;
      end
      8'h68 : begin
        _zz_io_ret = 8'h45;
      end
      8'h69 : begin
        _zz_io_ret = 8'hf9;
      end
      8'h6a : begin
        _zz_io_ret = 8'h02;
      end
      8'h6b : begin
        _zz_io_ret = 8'h7f;
      end
      8'h6c : begin
        _zz_io_ret = 8'h50;
      end
      8'h6d : begin
        _zz_io_ret = 8'h3c;
      end
      8'h6e : begin
        _zz_io_ret = 8'h9f;
      end
      8'h6f : begin
        _zz_io_ret = 8'ha8;
      end
      8'h70 : begin
        _zz_io_ret = 8'h51;
      end
      8'h71 : begin
        _zz_io_ret = 8'ha3;
      end
      8'h72 : begin
        _zz_io_ret = 8'h40;
      end
      8'h73 : begin
        _zz_io_ret = 8'h8f;
      end
      8'h74 : begin
        _zz_io_ret = 8'h92;
      end
      8'h75 : begin
        _zz_io_ret = 8'h9d;
      end
      8'h76 : begin
        _zz_io_ret = 8'h38;
      end
      8'h77 : begin
        _zz_io_ret = 8'hf5;
      end
      8'h78 : begin
        _zz_io_ret = 8'hbc;
      end
      8'h79 : begin
        _zz_io_ret = 8'hb6;
      end
      8'h7a : begin
        _zz_io_ret = 8'hda;
      end
      8'h7b : begin
        _zz_io_ret = 8'h21;
      end
      8'h7c : begin
        _zz_io_ret = 8'h10;
      end
      8'h7d : begin
        _zz_io_ret = 8'hff;
      end
      8'h7e : begin
        _zz_io_ret = 8'hf3;
      end
      8'h7f : begin
        _zz_io_ret = 8'hd2;
      end
      8'h80 : begin
        _zz_io_ret = 8'hcd;
      end
      8'h81 : begin
        _zz_io_ret = 8'h0c;
      end
      8'h82 : begin
        _zz_io_ret = 8'h13;
      end
      8'h83 : begin
        _zz_io_ret = 8'hec;
      end
      8'h84 : begin
        _zz_io_ret = 8'h5f;
      end
      8'h85 : begin
        _zz_io_ret = 8'h97;
      end
      8'h86 : begin
        _zz_io_ret = 8'h44;
      end
      8'h87 : begin
        _zz_io_ret = 8'h17;
      end
      8'h88 : begin
        _zz_io_ret = 8'hc4;
      end
      8'h89 : begin
        _zz_io_ret = 8'ha7;
      end
      8'h8a : begin
        _zz_io_ret = 8'h7e;
      end
      8'h8b : begin
        _zz_io_ret = 8'h3d;
      end
      8'h8c : begin
        _zz_io_ret = 8'h64;
      end
      8'h8d : begin
        _zz_io_ret = 8'h5d;
      end
      8'h8e : begin
        _zz_io_ret = 8'h19;
      end
      8'h8f : begin
        _zz_io_ret = 8'h73;
      end
      8'h90 : begin
        _zz_io_ret = 8'h60;
      end
      8'h91 : begin
        _zz_io_ret = 8'h81;
      end
      8'h92 : begin
        _zz_io_ret = 8'h4f;
      end
      8'h93 : begin
        _zz_io_ret = 8'hdc;
      end
      8'h94 : begin
        _zz_io_ret = 8'h22;
      end
      8'h95 : begin
        _zz_io_ret = 8'h2a;
      end
      8'h96 : begin
        _zz_io_ret = 8'h90;
      end
      8'h97 : begin
        _zz_io_ret = 8'h88;
      end
      8'h98 : begin
        _zz_io_ret = 8'h46;
      end
      8'h99 : begin
        _zz_io_ret = 8'hee;
      end
      8'h9a : begin
        _zz_io_ret = 8'hb8;
      end
      8'h9b : begin
        _zz_io_ret = 8'h14;
      end
      8'h9c : begin
        _zz_io_ret = 8'hde;
      end
      8'h9d : begin
        _zz_io_ret = 8'h5e;
      end
      8'h9e : begin
        _zz_io_ret = 8'h0b;
      end
      8'h9f : begin
        _zz_io_ret = 8'hdb;
      end
      8'ha0 : begin
        _zz_io_ret = 8'he0;
      end
      8'ha1 : begin
        _zz_io_ret = 8'h32;
      end
      8'ha2 : begin
        _zz_io_ret = 8'h3a;
      end
      8'ha3 : begin
        _zz_io_ret = 8'h0a;
      end
      8'ha4 : begin
        _zz_io_ret = 8'h49;
      end
      8'ha5 : begin
        _zz_io_ret = 8'h06;
      end
      8'ha6 : begin
        _zz_io_ret = 8'h24;
      end
      8'ha7 : begin
        _zz_io_ret = 8'h5c;
      end
      8'ha8 : begin
        _zz_io_ret = 8'hc2;
      end
      8'ha9 : begin
        _zz_io_ret = 8'hd3;
      end
      8'haa : begin
        _zz_io_ret = 8'hac;
      end
      8'hab : begin
        _zz_io_ret = 8'h62;
      end
      8'hac : begin
        _zz_io_ret = 8'h91;
      end
      8'had : begin
        _zz_io_ret = 8'h95;
      end
      8'hae : begin
        _zz_io_ret = 8'he4;
      end
      8'haf : begin
        _zz_io_ret = 8'h79;
      end
      8'hb0 : begin
        _zz_io_ret = 8'he7;
      end
      8'hb1 : begin
        _zz_io_ret = 8'hc8;
      end
      8'hb2 : begin
        _zz_io_ret = 8'h37;
      end
      8'hb3 : begin
        _zz_io_ret = 8'h6d;
      end
      8'hb4 : begin
        _zz_io_ret = 8'h8d;
      end
      8'hb5 : begin
        _zz_io_ret = 8'hd5;
      end
      8'hb6 : begin
        _zz_io_ret = 8'h4e;
      end
      8'hb7 : begin
        _zz_io_ret = 8'ha9;
      end
      8'hb8 : begin
        _zz_io_ret = 8'h6c;
      end
      8'hb9 : begin
        _zz_io_ret = 8'h56;
      end
      8'hba : begin
        _zz_io_ret = 8'hf4;
      end
      8'hbb : begin
        _zz_io_ret = 8'hea;
      end
      8'hbc : begin
        _zz_io_ret = 8'h65;
      end
      8'hbd : begin
        _zz_io_ret = 8'h7a;
      end
      8'hbe : begin
        _zz_io_ret = 8'hae;
      end
      8'hbf : begin
        _zz_io_ret = 8'h08;
      end
      8'hc0 : begin
        _zz_io_ret = 8'hba;
      end
      8'hc1 : begin
        _zz_io_ret = 8'h78;
      end
      8'hc2 : begin
        _zz_io_ret = 8'h25;
      end
      8'hc3 : begin
        _zz_io_ret = 8'h2e;
      end
      8'hc4 : begin
        _zz_io_ret = 8'h1c;
      end
      8'hc5 : begin
        _zz_io_ret = 8'ha6;
      end
      8'hc6 : begin
        _zz_io_ret = 8'hb4;
      end
      8'hc7 : begin
        _zz_io_ret = 8'hc6;
      end
      8'hc8 : begin
        _zz_io_ret = 8'he8;
      end
      8'hc9 : begin
        _zz_io_ret = 8'hdd;
      end
      8'hca : begin
        _zz_io_ret = 8'h74;
      end
      8'hcb : begin
        _zz_io_ret = 8'h1f;
      end
      8'hcc : begin
        _zz_io_ret = 8'h4b;
      end
      8'hcd : begin
        _zz_io_ret = 8'hbd;
      end
      8'hce : begin
        _zz_io_ret = 8'h8b;
      end
      8'hcf : begin
        _zz_io_ret = 8'h8a;
      end
      8'hd0 : begin
        _zz_io_ret = 8'h70;
      end
      8'hd1 : begin
        _zz_io_ret = 8'h3e;
      end
      8'hd2 : begin
        _zz_io_ret = 8'hb5;
      end
      8'hd3 : begin
        _zz_io_ret = 8'h66;
      end
      8'hd4 : begin
        _zz_io_ret = 8'h48;
      end
      8'hd5 : begin
        _zz_io_ret = 8'h03;
      end
      8'hd6 : begin
        _zz_io_ret = 8'hf6;
      end
      8'hd7 : begin
        _zz_io_ret = 8'h0e;
      end
      8'hd8 : begin
        _zz_io_ret = 8'h61;
      end
      8'hd9 : begin
        _zz_io_ret = 8'h35;
      end
      8'hda : begin
        _zz_io_ret = 8'h57;
      end
      8'hdb : begin
        _zz_io_ret = 8'hb9;
      end
      8'hdc : begin
        _zz_io_ret = 8'h86;
      end
      8'hdd : begin
        _zz_io_ret = 8'hc1;
      end
      8'hde : begin
        _zz_io_ret = 8'h1d;
      end
      8'hdf : begin
        _zz_io_ret = 8'h9e;
      end
      8'he0 : begin
        _zz_io_ret = 8'he1;
      end
      8'he1 : begin
        _zz_io_ret = 8'hf8;
      end
      8'he2 : begin
        _zz_io_ret = 8'h98;
      end
      8'he3 : begin
        _zz_io_ret = 8'h11;
      end
      8'he4 : begin
        _zz_io_ret = 8'h69;
      end
      8'he5 : begin
        _zz_io_ret = 8'hd9;
      end
      8'he6 : begin
        _zz_io_ret = 8'h8e;
      end
      8'he7 : begin
        _zz_io_ret = 8'h94;
      end
      8'he8 : begin
        _zz_io_ret = 8'h9b;
      end
      8'he9 : begin
        _zz_io_ret = 8'h1e;
      end
      8'hea : begin
        _zz_io_ret = 8'h87;
      end
      8'heb : begin
        _zz_io_ret = 8'he9;
      end
      8'hec : begin
        _zz_io_ret = 8'hce;
      end
      8'hed : begin
        _zz_io_ret = 8'h55;
      end
      8'hee : begin
        _zz_io_ret = 8'h28;
      end
      8'hef : begin
        _zz_io_ret = 8'hdf;
      end
      8'hf0 : begin
        _zz_io_ret = 8'h8c;
      end
      8'hf1 : begin
        _zz_io_ret = 8'ha1;
      end
      8'hf2 : begin
        _zz_io_ret = 8'h89;
      end
      8'hf3 : begin
        _zz_io_ret = 8'h0d;
      end
      8'hf4 : begin
        _zz_io_ret = 8'hbf;
      end
      8'hf5 : begin
        _zz_io_ret = 8'he6;
      end
      8'hf6 : begin
        _zz_io_ret = 8'h42;
      end
      8'hf7 : begin
        _zz_io_ret = 8'h68;
      end
      8'hf8 : begin
        _zz_io_ret = 8'h41;
      end
      8'hf9 : begin
        _zz_io_ret = 8'h99;
      end
      8'hfa : begin
        _zz_io_ret = 8'h2d;
      end
      8'hfb : begin
        _zz_io_ret = 8'h0f;
      end
      8'hfc : begin
        _zz_io_ret = 8'hb0;
      end
      8'hfd : begin
        _zz_io_ret = 8'h54;
      end
      8'hfe : begin
        _zz_io_ret = 8'hbb;
      end
      default : begin
        _zz_io_ret = 8'h16;
      end
    endcase
  end

  assign io_ret = _zz_io_ret;

endmodule
